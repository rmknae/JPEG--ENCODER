// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
//   Defines the standard 8x8 Discrete Cosine Transform (DCT) basis // matrix used in JPEG encoding and decoding.
//   - The matrix elements are based on the definition of the DCT-II.
//   - In hardware, these coefficients are usually scaled to fixed-point
//     representation (e.g., multiplied by 4096) 
//   - This version provides a fixed-point integer version (scaled by //4096), suitable for use in testbenches and hardware modules.
//
// Author : Rameen
// Date   : 29th July 2025
//


`ifndef DCT_CONSTANTS_SVH
`define DCT_CONSTANTS_SVH

`endif // DCT_CONSTANTS_SVH
