// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
//    Header file defining localparams for JPEG Huffman encoding.
//    - DC Huffman code lengths and codes (Luma & Chroma)
//    - AC Huffman code lengths and codes (Luma & Chroma)
//    - Run-length/size to Huffman index mapping
//
// Author: Rameen
// Date  : 23rd July 2025

`ifndef Y_HUFF_CONSTANTS_SVH
`define Y_HUFF_CONSTANTS_SVH

// -------------------- DC Code Lengths --------------------
parameter int Y_DC_code_length[0:11] = '{2,2,2,3,4,5,6,7,8,9,10,11};

// -------------------- DC Codes --------------------
parameter logic [10:0] Y_DC[0:11] = '{
    11'b00000000000, 11'b01000000000, 11'b10000000000, 11'b11000000000,
    11'b11100000000, 11'b11110000000, 11'b11111000000, 11'b11111100000,
    11'b11111110000, 11'b11111111000, 11'b11111111100, 11'b11111111110
};

// -------------------- AC Code Lengths --------------------
parameter int Y_AC_code_length[0:161] = '{
    2,2,3,4,4,4,5,5,5,6,6,7,7,7,7,8,
    8,8,9,9,9,9,9,10,10,10,10,10,11,11,11,11,
    12,12,12,12,15,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16
};

// -------------------- AC Codes --------------------
parameter logic [15:0] Y_AC[0:161] = '{
    16'b0000000000000000, 16'b0100000000000000, 16'b1000000000000000, 16'b1010000000000000,
    16'b1011000000000000, 16'b1100000000000000, 16'b1101000000000000, 16'b1101100000000000,
    16'b1110000000000000, 16'b1110100000000000, 16'b1110110000000000, 16'b1111000000000000,
    16'b1111001000000000, 16'b1111010000000000, 16'b1111011000000000, 16'b1111100000000000,
    16'b1111100100000000, 16'b1111101000000000, 16'b1111101100000000, 16'b1111101110000000,
    16'b1111110000000000, 16'b1111110010000000, 16'b1111110100000000, 16'b1111110110000000,
    16'b1111110111000000, 16'b1111111000000000, 16'b1111111001000000, 16'b1111111010000000,
    16'b1111111011000000, 16'b1111111011100000, 16'b1111111100000000, 16'b1111111100100000,
    16'b1111111101000000, 16'b1111111101010000, 16'b1111111101100000, 16'b1111111101110000,
    16'b1111111110000000, 16'b1111111110000010, 16'b1111111110000011, 16'b1111111110000100,
    16'b1111111110000101, 16'b1111111110000110, 16'b1111111110000111, 16'b1111111110001000,
    16'b1111111110001001, 16'b1111111110001010, 16'b1111111110001011, 16'b1111111110001100,
    16'b1111111110001101, 16'b1111111110001110, 16'b1111111110001111, 16'b1111111110010000,
    16'b1111111110010001, 16'b1111111110010010, 16'b1111111110010011, 16'b1111111110010100,
    16'b1111111110010101, 16'b1111111110010110, 16'b1111111110010111, 16'b1111111110011000,
    16'b1111111110011001, 16'b1111111110011010, 16'b1111111110011011, 16'b1111111110011100,
    16'b1111111110011101, 16'b1111111110011110, 16'b1111111110011111, 16'b1111111110100000,
    16'b1111111110100001, 16'b1111111110100010, 16'b1111111110100011, 16'b1111111110100100,
    16'b1111111110100101, 16'b1111111110100110, 16'b1111111110100111, 16'b1111111110101000,
    16'b1111111110101001, 16'b1111111110101010, 16'b1111111110101011, 16'b1111111110101100,
    16'b1111111110101101, 16'b1111111110101110, 16'b1111111110101111, 16'b1111111110110000,
    16'b1111111110110001, 16'b1111111110110010, 16'b1111111110110011, 16'b1111111110110100,
    16'b1111111110110101, 16'b1111111110110110, 16'b1111111110110111, 16'b1111111110111000,
    16'b1111111110111001, 16'b1111111110111010, 16'b1111111110111011, 16'b1111111110111100,
    16'b1111111110111101, 16'b1111111110111110, 16'b1111111110111111, 16'b1111111111000000,
    16'b1111111111000001, 16'b1111111111000010, 16'b1111111111000011, 16'b1111111111000100,
    16'b1111111111000101, 16'b1111111111000110, 16'b1111111111000111, 16'b1111111111001000,
    16'b1111111111001001, 16'b1111111111001010, 16'b1111111111001011, 16'b1111111111001100,
    16'b1111111111001101, 16'b1111111111001110, 16'b1111111111001111, 16'b1111111111010000,
    16'b1111111111010001, 16'b1111111111010010, 16'b1111111111010011, 16'b1111111111010100,
    16'b1111111111010101, 16'b1111111111010110, 16'b1111111111010111, 16'b1111111111011000,
    16'b1111111111011001, 16'b1111111111011010, 16'b1111111111011011, 16'b1111111111011100,
    16'b1111111111011101, 16'b1111111111011110, 16'b1111111111011111, 16'b1111111111100000,
    16'b1111111111100001, 16'b1111111111100010, 16'b1111111111100011, 16'b1111111111100100,
    16'b1111111111100101, 16'b1111111111100110, 16'b1111111111100111, 16'b1111111111101000,
    16'b1111111111101001, 16'b1111111111101010, 16'b1111111111101011, 16'b1111111111101100,
    16'b1111111111101101, 16'b1111111111101110, 16'b1111111111101111, 16'b1111111111110000,
    16'b1111111111110001, 16'b1111111111110010, 16'b1111111111110011, 16'b1111111111110100,
    16'b1111111111110101, 16'b1111111111110110, 16'b1111111111110111, 16'b1111111111111000,
    16'b1111111111111001, 16'b1111111111111010, 16'b1111111111111011, 16'b1111111111111100,
    16'b1111111111111101, 16'b1111111111111110
};

parameter int Y_AC_run_code [0:250] = '{
        // Explicit assignments
        0: 3,  1: 0,  2: 1,  3: 2,  4: 4,
        5: 6,  6: 11, 7: 15, 8: 23, 9: 37,
        10: 38, 11: 0, 12: 0, 13: 0, 14: 0, 15: 0,
        16: 0, 17: 5, 18: 7, 19: 12, 20: 18,
        21: 28, 22: 39, 23: 40, 24: 41, 25: 42,
        26: 43, 27: 0, 28: 0, 29: 0, 30: 0, 31: 0,
        32: 0, 33: 8, 34: 16, 35: 24, 36: 32,
        37: 44, 38: 45, 39: 46, 40: 47, 41: 48,
        42: 49, 43: 0, 44: 0, 45: 0, 46: 0, 47: 0,
        48: 0, 49: 9, 50: 19, 51: 33, 52: 50,
        53: 51, 54: 52, 55: 53, 56: 54, 57: 55,
        58: 56, 59: 0, 60: 0, 61: 0, 62: 0, 63: 0,
        64: 0, 65: 10, 66: 25, 67: 57, 68: 58,
        69: 59, 70: 60, 71: 61, 72: 62, 73: 63,
        74: 64, 75: 0, 76: 0, 77: 0, 78: 0, 79: 0,
        80: 0, 81: 13, 82: 29, 83: 65, 84: 66,
        85: 67, 86: 68, 87: 69, 88: 70, 89: 71,
        90: 72, 91: 0, 92: 0, 93: 0, 94: 0, 95: 0,
        96: 0, 97: 14, 98: 34, 99: 73, 100: 74,
        101: 75, 102: 76, 103: 77, 104: 78, 105: 79,
        106: 80, 107: 0, 108: 0, 109: 0, 110: 0, 111: 0,
        112: 0, 113: 17, 114: 35, 115: 81, 116: 82,
        117: 83, 118: 84, 119: 85, 120: 86, 121: 87,
        122: 88, 123: 0, 124: 0, 125: 0, 126: 0, 127: 0,
        128: 0, 129: 20, 130: 36, 131: 89, 132: 90,
        133: 91, 134: 92, 135: 93, 136: 94, 137: 95,
        138: 96, 139: 0, 140: 0, 141: 0, 142: 0, 143: 0,
        144: 0, 145: 21, 146: 97, 147: 98, 148: 99,
        149: 100,150: 101,151: 102,152: 103,153: 104,
        154: 105,155: 0, 156: 0, 157: 0, 158: 0, 159: 0,
        160: 0, 161: 22, 162: 106,163: 107,164: 108,
        165: 109,166: 110,167: 111,168: 112,169: 113,
        170: 114,171: 0, 172: 0, 173: 0, 174: 0, 175: 0,
        176: 0, 177: 26, 178: 115,179: 116,180: 117,
        181: 118,182: 119,183: 120,184: 121,185: 122,
        186: 123,187: 0, 188: 0, 189: 0, 190: 0, 191: 0,
        192: 0, 193: 27, 194: 124,195: 125,196: 126,
        197: 127,198: 128,199: 129,200: 130,201: 131,
        202: 132,203: 0, 204: 0, 205: 0, 206: 0, 207: 0,
        208: 0, 209: 30, 210: 133,211: 134,212: 135,
        213: 136,214: 137,215: 138,216: 139,217: 140,
        218: 141,219: 0, 220: 0, 221: 0, 222: 0, 223: 0,
        224: 0, 225: 142,226: 143,227: 144,228: 145,
        229: 146,230: 147,231: 148,232: 149,233: 150,
        234: 151,235: 0, 236: 0, 237: 0, 238: 0, 239: 0,
        240: 31, 241: 152,242: 153,243: 154,244: 155,
        245: 156,246: 157,247: 158,248: 159,249: 160,
        250: 161,

        // Default fill for all unspecified = 0
        default: 0
    };
`endif //y_ HUFF_CONSTANTS_SVH
