		
`timescale 1ps/1ps

module jpeg_top_tb;

    // ----------------------
    // Declarations
    // ----------------------
    logic end_of_file_signal;
    logic [23:0] data_in;
    logic clk;
    logic rst;
    logic enable;
  logic yes;
    wire [31:0] JPEG_bitstream;
    wire data_ready;
    wire [4:0] end_of_file_bitstream_count;
    wire eof_data_partial_ready;

    integer outfile;

    // ----------------------
    // Unit Under Test
    // ----------------------
    jpeg_top UUT (
        .end_of_file_signal(end_of_file_signal),
        .data_in(data_in),
        .clk(clk),
        .rst(rst),
        .enable(enable),
        .JPEG_bitstream(JPEG_bitstream),
        .data_ready(data_ready),
        .end_of_file_bitstream_count(end_of_file_bitstream_count),
        .eof_data_partial_ready(eof_data_partial_ready)
    );

    // ----------------------
    // Stimulus process
    // ----------------------
    initial begin : STIMUL
        rst = 1'b1;
        enable = 1'b0;
        end_of_file_signal = 1'b0;
        data_in = '0;
   yes = 1'b0;
        #10000;
        rst = 1'b0;
        enable = 1'b1;

	
	
	data_in <= 24'b010100100011000100000101;
#10000;
	data_in <= 24'b010100100011000100000110;
#10000;
	data_in <= 24'b010100110011001100000110;
#10000;
	data_in <= 24'b010100110011001100000111;
#10000;
	data_in <= 24'b010101000011010000001000;
#10000;
	data_in <= 24'b010101010011010100001000;
#10000;
	data_in <= 24'b010101100011011000001001;
#10000;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010100110011001000000101;
#10000;
	data_in <= 24'b010101000011010000000110;
#10000;
	data_in <= 24'b010101000011010000000111;
#10000;
	data_in <= 24'b010101010011010100001000;
#10000;
	data_in <= 24'b010101010011010100001001;
#10000;
	data_in <= 24'b010101010011010100001010;
#10000;
	data_in <= 24'b010101100011010100001011;
#10000;
	data_in <= 24'b010101110011011100001100;
#10000;
	data_in <= 24'b010101010011010100000110;
#10000;
	data_in <= 24'b010101010011010100000111;
#10000;
	data_in <= 24'b010101100011011000001001;
#10000;
	data_in <= 24'b010101100011011000001001;
#10000;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010101110011011100001011;
#10000;
	data_in <= 24'b010101110011100000001100;
#10000;
	data_in <= 24'b010110000011101000001101;
#10000;
	data_in <= 24'b010101010011010100001001;
#10000;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010101110011011100001011;
#10000;
	data_in <= 24'b010110000011100000001101;
#10000;
	data_in <= 24'b010110000011100000001110;
#10000;
	data_in <= 24'b010110010011100100001110;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b010101100011011100001011;
#10000;
	data_in <= 24'b010101110011011100001011;
#10000;
	data_in <= 24'b010110000011100000001100;
#10000;
	data_in <= 24'b010110000011100100001110;
#10000;
	data_in <= 24'b010110000011101000001101;
#10000;
	data_in <= 24'b010110010011101100001110;
#10000;
	data_in <= 24'b010110110011101100001111;
#10000;
	data_in <= 24'b010111000011110000010001;
#10000;
	data_in <= 24'b010110000011100000001011;
#10000;
	data_in <= 24'b010110000011100100001100;
#10000;
	data_in <= 24'b010110010011101000001110;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b010110100011110000001111;
#10000;
	data_in <= 24'b010110110011110100001111;
#10000;
	data_in <= 24'b010111000011110100010001;
#10000;
	data_in <= 24'b010111010011111000010010;
#10000;
	data_in <= 24'b010110000011100000001011;
#10000;
	data_in <= 24'b010110100011101000001101;
#10000;
	data_in <= 24'b010110100011101100001110;
#10000;
	data_in <= 24'b010110110011110100001111;
#10000;
	data_in <= 24'b010111000011110100010000;
#10000;
	data_in <= 24'b010111010011111000010001;
#10000;
	data_in <= 24'b010111100011111100010011;
#10000;
	data_in <= 24'b010111110100000000010100;
#10000;
	data_in <= 24'b010110100011101000001110;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b010110110011110100010000;
#10000;
	data_in <= 24'b010111010011111000010001;
#10000;
	data_in <= 24'b010111100011111100010010;
#10000;
	data_in <= 24'b010111110100000000010100;
#10000;
	data_in <= 24'b011000000100001000010101;
#10000;
	data_in <= 24'b011000010100001100010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010101100011011000001011;
#10000;
	data_in <= 24'b010101110011011100001100;
#10000;
	data_in <= 24'b010101110011100000001100;
#10000;
	data_in <= 24'b010101110011100000001100;
#10000;
	data_in <= 24'b010110000011100000001101;
#10000;
	data_in <= 24'b010110010011101000001111;
#10000;
	data_in <= 24'b010110010011101000001111;
#10000;
	data_in <= 24'b010110010011101000001111;
#10000;
	data_in <= 24'b010101110011100000001011;
#10000;
	data_in <= 24'b010110000011100100001101;
#10000;
	data_in <= 24'b010110010011101000001110;
#10000;
	data_in <= 24'b010110010011100100001110;
#10000;
	data_in <= 24'b010110100011101000001111;
#10000;
	data_in <= 24'b010110110011101100010000;
#10000;
	data_in <= 24'b010110100011101100010000;
#10000;
	data_in <= 24'b010110100011110000010001;
#10000;
	data_in <= 24'b010110010011101000001101;
#10000;
	data_in <= 24'b010110100011101000001110;
#10000;
	data_in <= 24'b010110110011101100001111;
#10000;
	data_in <= 24'b010110110011101100010000;
#10000;
	data_in <= 24'b010110110011110000010001;
#10000;
	data_in <= 24'b010111000011110100010010;
#10000;
	data_in <= 24'b010111000011110100010010;
#10000;
	data_in <= 24'b010111000011110100010010;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b010110110011101100010001;
#10000;
	data_in <= 24'b010111000011110100010001;
#10000;
	data_in <= 24'b010111000011110100010001;
#10000;
	data_in <= 24'b010111010011111000010011;
#10000;
	data_in <= 24'b010111010011111000010100;
#10000;
	data_in <= 24'b010111010011111000010100;
#10000;
	data_in <= 24'b010111100011111100010101;
#10000;
	data_in <= 24'b010110110011110000010010;
#10000;
	data_in <= 24'b010111010011111000010010;
#10000;
	data_in <= 24'b010111000011111100010011;
#10000;
	data_in <= 24'b010111010100000000010100;
#10000;
	data_in <= 24'b010111110100000000010101;
#10000;
	data_in <= 24'b010111110100000000010110;
#10000;
	data_in <= 24'b010111110100000100010111;
#10000;
	data_in <= 24'b011000000100001000011000;
#10000;
	data_in <= 24'b010111010011111100010011;
#10000;
	data_in <= 24'b010111100100000000010100;
#10000;
	data_in <= 24'b010111110100000100010110;
#10000;
	data_in <= 24'b010111110100001100010110;
#10000;
	data_in <= 24'b011000000100001100010111;
#10000;
	data_in <= 24'b011000010100001100011000;
#10000;
	data_in <= 24'b011000100100001100011010;
#10000;
	data_in <= 24'b011000100100010000011010;
#10000;
	data_in <= 24'b010111110100000100010100;
#10000;
	data_in <= 24'b011000000100001000010110;
#10000;
	data_in <= 24'b011000000100001100010111;
#10000;
	data_in <= 24'b011000010100010000011000;
#10000;
	data_in <= 24'b011000010100010000011001;
#10000;
	data_in <= 24'b011000100100010100011010;
#10000;
	data_in <= 24'b011000110100011000011011;
#10000;
	data_in <= 24'b011001000100011100011100;
#10000;
	data_in <= 24'b011000010100001100011000;
#10000;
	data_in <= 24'b011000100100010000011000;
#10000;
	data_in <= 24'b011000100100010000011001;
#10000;
	data_in <= 24'b011000100100010000011011;
#10000;
	data_in <= 24'b011000110100011000011100;
#10000;
	data_in <= 24'b011001000100100000011100;
#10000;
	data_in <= 24'b011001000100100000011101;
#10000;
	data_in <= 24'b011001100100100000011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010110010011101100010000;
#10000;
	data_in <= 24'b010110100011110000010001;
#10000;
	data_in <= 24'b010110100011110000010010;
#10000;
	data_in <= 24'b010110100011110000010010;
#10000;
	data_in <= 24'b010110100011110000010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010011;
#10000;
	data_in <= 24'b010110110011111000010100;
#10000;
	data_in <= 24'b010111000011111000010100;
#10000;
	data_in <= 24'b010111010100000000010101;
#10000;
	data_in <= 24'b010111100100000000010101;
#10000;
	data_in <= 24'b010111010011111000010011;
#10000;
	data_in <= 24'b010111010011111100010100;
#10000;
	data_in <= 24'b010111010011111100010100;
#10000;
	data_in <= 24'b010111010100000000010101;
#10000;
	data_in <= 24'b010111100100000100010110;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100001000010111;
#10000;
	data_in <= 24'b010111110100001000010111;
#10000;
	data_in <= 24'b010111100011111100010101;
#10000;
	data_in <= 24'b010111100100000100010110;
#10000;
	data_in <= 24'b010111110100001000011000;
#10000;
	data_in <= 24'b010111110100001000011000;
#10000;
	data_in <= 24'b011000000100001100011000;
#10000;
	data_in <= 24'b011000000100001100011001;
#10000;
	data_in <= 24'b011000000100001100011010;
#10000;
	data_in <= 24'b011000010100010000011011;
#10000;
	data_in <= 24'b011000010100001100011000;
#10000;
	data_in <= 24'b011000000100001100011001;
#10000;
	data_in <= 24'b011000010100010000011010;
#10000;
	data_in <= 24'b011000100100010100011011;
#10000;
	data_in <= 24'b011000010100010100011011;
#10000;
	data_in <= 24'b011000100100011000011100;
#10000;
	data_in <= 24'b011000110100010100011100;
#10000;
	data_in <= 24'b011000110100011000011101;
#10000;
	data_in <= 24'b011000100100010100011010;
#10000;
	data_in <= 24'b011000110100011100011011;
#10000;
	data_in <= 24'b011000110100011100011100;
#10000;
	data_in <= 24'b011000110100011100011101;
#10000;
	data_in <= 24'b011001000100100000011110;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001100100100100100000;
#10000;
	data_in <= 24'b011001000100011100011100;
#10000;
	data_in <= 24'b011001010100100000011101;
#10000;
	data_in <= 24'b011001010100100100011110;
#10000;
	data_in <= 24'b011001100100100100011110;
#10000;
	data_in <= 24'b011001100100101000100000;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100100100100000;
#10000;
	data_in <= 24'b011010000100101000100000;
#10000;
	data_in <= 24'b011010000100101100100001;
#10000;
	data_in <= 24'b011010010100110100100011;
#10000;
	data_in <= 24'b011010010100110100100100;
#10000;
	data_in <= 24'b011010100100111000100100;
#10000;
	data_in <= 24'b011010100100111000100100;
#10000;
	data_in <= 24'b011010100100111000100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111000011111000010100;
#10000;
	data_in <= 24'b010111000011111000010100;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111010100000000010101;
#10000;
	data_in <= 24'b010111010100000100010110;
#10000;
	data_in <= 24'b010111010100000000010110;
#10000;
	data_in <= 24'b010111100100000100010110;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100000100011000;
#10000;
	data_in <= 24'b011000000100001100011000;
#10000;
	data_in <= 24'b011000000100001100011000;
#10000;
	data_in <= 24'b011000000100001100011001;
#10000;
	data_in <= 24'b011000000100001100011010;
#10000;
	data_in <= 24'b011000010100001100011010;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100010000011011;
#10000;
	data_in <= 24'b011000100100010000011011;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011001000100011000011110;
#10000;
	data_in <= 24'b011001000100011100011110;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100100100001;
#10000;
	data_in <= 24'b011001100100101000100001;
#10000;
	data_in <= 24'b011001100100101000100001;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100101100100010;
#10000;
	data_in <= 24'b011001110100110000100011;
#10000;
	data_in <= 24'b011010000100110000100011;
#10000;
	data_in <= 24'b011010000100110000100011;
#10000;
	data_in <= 24'b011010000100110000100010;
#10000;
	data_in <= 24'b011010010100110100100011;
#10000;
	data_in <= 24'b011010010100110100100011;
#10000;
	data_in <= 24'b011010010100110100100100;
#10000;
	data_in <= 24'b011010010100111000100101;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010100100111100100110;
#10000;
	data_in <= 24'b011010100100111100100110;
#10000;
	data_in <= 24'b011010100100111100100110;
#10000;
	data_in <= 24'b011010110100111100100111;
#10000;
	data_in <= 24'b011010110101000000101000;
#10000;
	data_in <= 24'b011011000101000100101000;
#10000;
	data_in <= 24'b011011000101000100101000;
#10000;
	data_in <= 24'b011011000101000100101001;
#10000;
	data_in <= 24'b011011010101001000101010;
#10000;
	data_in <= 24'b011011000101001000101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111000100000000010110;
#10000;
	data_in <= 24'b010111000100000000010110;
#10000;
	data_in <= 24'b010111000100000000010111;
#10000;
	data_in <= 24'b010111000100000000010111;
#10000;
	data_in <= 24'b010111010100000000011000;
#10000;
	data_in <= 24'b010111010100000000011001;
#10000;
	data_in <= 24'b010111010100000000011000;
#10000;
	data_in <= 24'b010111010100000000011000;
#10000;
	data_in <= 24'b010111100100000100011000;
#10000;
	data_in <= 24'b010111110100001000011001;
#10000;
	data_in <= 24'b010111110100001100011010;
#10000;
	data_in <= 24'b010111110100001000011001;
#10000;
	data_in <= 24'b010111110100001000011001;
#10000;
	data_in <= 24'b011000000100001000011010;
#10000;
	data_in <= 24'b011000000100001000011010;
#10000;
	data_in <= 24'b011000000100001100011011;
#10000;
	data_in <= 24'b011000010100010000011011;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011101;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011100011110;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011001000100011100100000;
#10000;
	data_in <= 24'b011001000100011100100000;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001010100100100100001;
#10000;
	data_in <= 24'b011001010100100100100001;
#10000;
	data_in <= 24'b011001010100100100100010;
#10000;
	data_in <= 24'b011001010100101000100010;
#10000;
	data_in <= 24'b011001100100101000100010;
#10000;
	data_in <= 24'b011001010100101100100010;
#10000;
	data_in <= 24'b011001100100101000100011;
#10000;
	data_in <= 24'b011001110100101000100100;
#10000;
	data_in <= 24'b011010000100110000100100;
#10000;
	data_in <= 24'b011010000100110000100101;
#10000;
	data_in <= 24'b011010000100110100100101;
#10000;
	data_in <= 24'b011010000100110100100101;
#10000;
	data_in <= 24'b011010000100111000100101;
#10000;
	data_in <= 24'b011010000100111000100101;
#10000;
	data_in <= 24'b011010000100111000100101;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010100100111100100111;
#10000;
	data_in <= 24'b011010100100111100101000;
#10000;
	data_in <= 24'b011010100100111100100111;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011011010101001000101011;
#10000;
	data_in <= 24'b011011010101001000101100;
#10000;
	data_in <= 24'b011011010101001000101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011110101001100101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111100100000000011000;
#10000;
	data_in <= 24'b010111100100000000011000;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001000100100000100001;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001100100101000100100;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100101000100011;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100110000100101;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010010100111000100111;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011011110101001100101101;
#10000;
	data_in <= 24'b011011110101001100101101;
#10000;
	data_in <= 24'b011011110101001100101100;
#10000;
	data_in <= 24'b011011110101001100101101;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101110;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000100011001;
#10000;
	data_in <= 24'b010111100100000000011000;
#10000;
	data_in <= 24'b010111100100000000011000;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100010000011100;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001000100100000100010;
#10000;
	data_in <= 24'b011001000100100000100001;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100110000100101;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100101000100011;
#10000;
	data_in <= 24'b011001100100101100100100;
#10000;
	data_in <= 24'b011001100100101000100100;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010010100111100100111;
#10000;
	data_in <= 24'b011010010100111000100111;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000100101010;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011011110101010000101110;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101110;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101001100101101;
#10000;
	data_in <= 24'b011011110101001100101100;
#10000;
	data_in <= 24'b011011110101001100101101;
#10000;
	data_in <= 24'b011011110101001100101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111010100000000011000;
#10000;
	data_in <= 24'b010111010100000000011000;
#10000;
	data_in <= 24'b010111010100000000011001;
#10000;
	data_in <= 24'b010111010100000000011000;
#10000;
	data_in <= 24'b010111000100000000010111;
#10000;
	data_in <= 24'b010111000100000000010111;
#10000;
	data_in <= 24'b010111000100000000010110;
#10000;
	data_in <= 24'b010111000100000000010110;
#10000;
	data_in <= 24'b011000000100001100011011;
#10000;
	data_in <= 24'b011000000100001000011010;
#10000;
	data_in <= 24'b011000000100001000011010;
#10000;
	data_in <= 24'b010111110100001000011001;
#10000;
	data_in <= 24'b010111110100001000011001;
#10000;
	data_in <= 24'b010111110100001100011010;
#10000;
	data_in <= 24'b010111110100001000011001;
#10000;
	data_in <= 24'b010111100100000100011000;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000100100010100011101;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000010100010000011011;
#10000;
	data_in <= 24'b011001000100011100100001;
#10000;
	data_in <= 24'b011001000100011100100000;
#10000;
	data_in <= 24'b011001000100011100100000;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011111;
#10000;
	data_in <= 24'b011000110100011100011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011001110100101000100100;
#10000;
	data_in <= 24'b011001100100101000100011;
#10000;
	data_in <= 24'b011001010100101100100010;
#10000;
	data_in <= 24'b011001100100101000100010;
#10000;
	data_in <= 24'b011001010100101000100010;
#10000;
	data_in <= 24'b011001010100100100100010;
#10000;
	data_in <= 24'b011001010100100100100001;
#10000;
	data_in <= 24'b011001010100100100100001;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010000100111000100101;
#10000;
	data_in <= 24'b011010000100111000100101;
#10000;
	data_in <= 24'b011010000100111000100101;
#10000;
	data_in <= 24'b011010000100110100100101;
#10000;
	data_in <= 24'b011010000100110100100101;
#10000;
	data_in <= 24'b011010000100110000100101;
#10000;
	data_in <= 24'b011010000100110000100100;
#10000;
	data_in <= 24'b011010110101000000101001;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010100101000000101000;
#10000;
	data_in <= 24'b011010100100111100100111;
#10000;
	data_in <= 24'b011010100100111100101000;
#10000;
	data_in <= 24'b011010100100111100100111;
#10000;
	data_in <= 24'b011011110101001100101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011010101001100101100;
#10000;
	data_in <= 24'b011011010101001000101100;
#10000;
	data_in <= 24'b011011010101001000101100;
#10000;
	data_in <= 24'b011011010101001000101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111100010101;
#10000;
	data_in <= 24'b010111000011111000010100;
#10000;
	data_in <= 24'b010111000011111000010100;
#10000;
	data_in <= 24'b010111100100000100011000;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100000100010110;
#10000;
	data_in <= 24'b010111010100000000010110;
#10000;
	data_in <= 24'b010111010100000100010110;
#10000;
	data_in <= 24'b010111010100000000010101;
#10000;
	data_in <= 24'b011000010100010000011011;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100001100011011;
#10000;
	data_in <= 24'b011000010100001100011010;
#10000;
	data_in <= 24'b011000000100001100011010;
#10000;
	data_in <= 24'b011000000100001100011001;
#10000;
	data_in <= 24'b011000000100001100011000;
#10000;
	data_in <= 24'b011000000100001100011000;
#10000;
	data_in <= 24'b011001000100011000011110;
#10000;
	data_in <= 24'b011000110100011000011110;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000110100010100011101;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010100011100;
#10000;
	data_in <= 24'b011000100100010000011011;
#10000;
	data_in <= 24'b011001010100100100100001;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100100100000;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001000100011100011110;
#10000;
	data_in <= 24'b011010000100110000100011;
#10000;
	data_in <= 24'b011010000100110000100011;
#10000;
	data_in <= 24'b011001110100110000100011;
#10000;
	data_in <= 24'b011001110100101100100010;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001100100101000100001;
#10000;
	data_in <= 24'b011001100100101000100001;
#10000;
	data_in <= 24'b011010100100111100100110;
#10000;
	data_in <= 24'b011010100100111100100110;
#10000;
	data_in <= 24'b011010010100111000100110;
#10000;
	data_in <= 24'b011010010100111000100101;
#10000;
	data_in <= 24'b011010010100110100100100;
#10000;
	data_in <= 24'b011010010100110100100011;
#10000;
	data_in <= 24'b011010010100110100100011;
#10000;
	data_in <= 24'b011010000100110000100010;
#10000;
	data_in <= 24'b011011000101001000101011;
#10000;
	data_in <= 24'b011011010101001000101010;
#10000;
	data_in <= 24'b011011000101000100101001;
#10000;
	data_in <= 24'b011011000101000100101000;
#10000;
	data_in <= 24'b011011000101000100101000;
#10000;
	data_in <= 24'b011010110101000000101000;
#10000;
	data_in <= 24'b011010110100111100100111;
#10000;
	data_in <= 24'b011010100100111100100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110100011110000010010;
#10000;
	data_in <= 24'b010110100011110000010010;
#10000;
	data_in <= 24'b010110100011110000010010;
#10000;
	data_in <= 24'b010110100011110000010001;
#10000;
	data_in <= 24'b010110010011101100010000;
#10000;
	data_in <= 24'b010111100100000000010101;
#10000;
	data_in <= 24'b010111010100000000010101;
#10000;
	data_in <= 24'b010111000011111000010100;
#10000;
	data_in <= 24'b010110110011111000010100;
#10000;
	data_in <= 24'b010110110011110100010011;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010110110011110100010010;
#10000;
	data_in <= 24'b010111110100001000010111;
#10000;
	data_in <= 24'b010111100100001000010111;
#10000;
	data_in <= 24'b010111100100000100010111;
#10000;
	data_in <= 24'b010111100100000100010110;
#10000;
	data_in <= 24'b010111010100000000010101;
#10000;
	data_in <= 24'b010111010011111100010100;
#10000;
	data_in <= 24'b010111010011111100010100;
#10000;
	data_in <= 24'b010111010011111000010011;
#10000;
	data_in <= 24'b011000010100010000011011;
#10000;
	data_in <= 24'b011000000100001100011010;
#10000;
	data_in <= 24'b011000000100001100011001;
#10000;
	data_in <= 24'b011000000100001100011000;
#10000;
	data_in <= 24'b010111110100001000011000;
#10000;
	data_in <= 24'b010111110100001000011000;
#10000;
	data_in <= 24'b010111100100000100010110;
#10000;
	data_in <= 24'b010111100011111100010101;
#10000;
	data_in <= 24'b011000110100011000011101;
#10000;
	data_in <= 24'b011000110100010100011100;
#10000;
	data_in <= 24'b011000100100011000011100;
#10000;
	data_in <= 24'b011000010100010100011011;
#10000;
	data_in <= 24'b011000100100010100011011;
#10000;
	data_in <= 24'b011000010100010000011010;
#10000;
	data_in <= 24'b011000000100001100011001;
#10000;
	data_in <= 24'b011000010100001100011000;
#10000;
	data_in <= 24'b011001100100100100100000;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001000100100000011110;
#10000;
	data_in <= 24'b011000110100011100011101;
#10000;
	data_in <= 24'b011000110100011100011100;
#10000;
	data_in <= 24'b011000110100011100011011;
#10000;
	data_in <= 24'b011000100100010100011010;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001100100101000100000;
#10000;
	data_in <= 24'b011001100100100100011110;
#10000;
	data_in <= 24'b011001010100100100011110;
#10000;
	data_in <= 24'b011001010100100000011101;
#10000;
	data_in <= 24'b011001000100011100011100;
#10000;
	data_in <= 24'b011010100100111000100101;
#10000;
	data_in <= 24'b011010100100111000100100;
#10000;
	data_in <= 24'b011010100100111000100100;
#10000;
	data_in <= 24'b011010010100110100100100;
#10000;
	data_in <= 24'b011010010100110100100011;
#10000;
	data_in <= 24'b011010000100101100100001;
#10000;
	data_in <= 24'b011010000100101000100000;
#10000;
	data_in <= 24'b011001110100100100100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010110010011101000001111;
#10000;
	data_in <= 24'b010110010011101000001111;
#10000;
	data_in <= 24'b010110010011101000001111;
#10000;
	data_in <= 24'b010110000011100000001101;
#10000;
	data_in <= 24'b010101110011100000001100;
#10000;
	data_in <= 24'b010101110011100000001100;
#10000;
	data_in <= 24'b010101110011011100001100;
#10000;
	data_in <= 24'b010101100011011000001011;
#10000;
	data_in <= 24'b010110100011110000010001;
#10000;
	data_in <= 24'b010110100011101100010000;
#10000;
	data_in <= 24'b010110110011101100010000;
#10000;
	data_in <= 24'b010110100011101000001111;
#10000;
	data_in <= 24'b010110010011100100001110;
#10000;
	data_in <= 24'b010110010011101000001110;
#10000;
	data_in <= 24'b010110000011100100001101;
#10000;
	data_in <= 24'b010101110011100000001011;
#10000;
	data_in <= 24'b010111000011110100010010;
#10000;
	data_in <= 24'b010111000011110100010010;
#10000;
	data_in <= 24'b010111000011110100010010;
#10000;
	data_in <= 24'b010110110011110000010001;
#10000;
	data_in <= 24'b010110110011101100010000;
#10000;
	data_in <= 24'b010110110011101100001111;
#10000;
	data_in <= 24'b010110100011101000001110;
#10000;
	data_in <= 24'b010110010011101000001101;
#10000;
	data_in <= 24'b010111100011111100010101;
#10000;
	data_in <= 24'b010111010011111000010100;
#10000;
	data_in <= 24'b010111010011111000010100;
#10000;
	data_in <= 24'b010111010011111000010011;
#10000;
	data_in <= 24'b010111000011110100010001;
#10000;
	data_in <= 24'b010111000011110100010001;
#10000;
	data_in <= 24'b010110110011101100010001;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b011000000100001000011000;
#10000;
	data_in <= 24'b010111110100000100010111;
#10000;
	data_in <= 24'b010111110100000000010110;
#10000;
	data_in <= 24'b010111110100000000010101;
#10000;
	data_in <= 24'b010111010100000000010100;
#10000;
	data_in <= 24'b010111000011111100010011;
#10000;
	data_in <= 24'b010111010011111000010010;
#10000;
	data_in <= 24'b010110110011110000010010;
#10000;
	data_in <= 24'b011000100100010000011010;
#10000;
	data_in <= 24'b011000100100001100011010;
#10000;
	data_in <= 24'b011000010100001100011000;
#10000;
	data_in <= 24'b011000000100001100010111;
#10000;
	data_in <= 24'b010111110100001100010110;
#10000;
	data_in <= 24'b010111110100000100010110;
#10000;
	data_in <= 24'b010111100100000000010100;
#10000;
	data_in <= 24'b010111010011111100010011;
#10000;
	data_in <= 24'b011001000100011100011100;
#10000;
	data_in <= 24'b011000110100011000011011;
#10000;
	data_in <= 24'b011000100100010100011010;
#10000;
	data_in <= 24'b011000010100010000011001;
#10000;
	data_in <= 24'b011000010100010000011000;
#10000;
	data_in <= 24'b011000000100001100010111;
#10000;
	data_in <= 24'b011000000100001000010110;
#10000;
	data_in <= 24'b010111110100000100010100;
#10000;
	data_in <= 24'b011001100100100000011111;
#10000;
	data_in <= 24'b011001000100100000011101;
#10000;
	data_in <= 24'b011001000100100000011100;
#10000;
	data_in <= 24'b011000110100011000011100;
#10000;
	data_in <= 24'b011000100100010000011011;
#10000;
	data_in <= 24'b011000100100010000011001;
#10000;
	data_in <= 24'b011000100100010000011000;
#10000;
	data_in <= 24'b011000010100001100011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010101100011011000001001;
#10000;
	data_in <= 24'b010101010011010100001000;
#10000;
	data_in <= 24'b010101000011010000001000;
#10000;
	data_in <= 24'b010100110011001100000111;
#10000;
	data_in <= 24'b010100110011001100000110;
#10000;
	data_in <= 24'b010100100011000100000110;
#10000;
	data_in <= 24'b010100100011000100000101;
#10000;
	data_in <= 24'b010101110011011100001100;
#10000;
	data_in <= 24'b010101100011010100001011;
#10000;
	data_in <= 24'b010101010011010100001010;
#10000;
	data_in <= 24'b010101010011010100001001;
#10000;
	data_in <= 24'b010101010011010100001000;
#10000;
	data_in <= 24'b010101000011010000000111;
#10000;
	data_in <= 24'b010101000011010000000110;
#10000;
	data_in <= 24'b010100110011001000000101;
#10000;
	data_in <= 24'b010110000011101000001101;
#10000;
	data_in <= 24'b010101110011100000001100;
#10000;
	data_in <= 24'b010101110011011100001011;
#10000;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010101100011011000001001;
#10000;
	data_in <= 24'b010101100011011000001001;
#10000;
	data_in <= 24'b010101010011010100000111;
#10000;
	data_in <= 24'b010101010011010100000110;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b010110010011100100001110;
#10000;
	data_in <= 24'b010110000011100000001110;
#10000;
	data_in <= 24'b010110000011100000001101;
#10000;
	data_in <= 24'b010101110011011100001011;
#10000;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010101100011011000001010;
#10000;
	data_in <= 24'b010101010011010100001001;
#10000;
	data_in <= 24'b010111000011110000010001;
#10000;
	data_in <= 24'b010110110011101100001111;
#10000;
	data_in <= 24'b010110010011101100001110;
#10000;
	data_in <= 24'b010110000011101000001101;
#10000;
	data_in <= 24'b010110000011100100001110;
#10000;
	data_in <= 24'b010110000011100000001100;
#10000;
	data_in <= 24'b010101110011011100001011;
#10000;
	data_in <= 24'b010101100011011100001011;
#10000;
	data_in <= 24'b010111010011111000010010;
#10000;
	data_in <= 24'b010111000011110100010001;
#10000;
	data_in <= 24'b010110110011110100001111;
#10000;
	data_in <= 24'b010110100011110000001111;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b010110010011101000001110;
#10000;
	data_in <= 24'b010110000011100100001100;
#10000;
	data_in <= 24'b010110000011100000001011;
#10000;
	data_in <= 24'b010111110100000000010100;
#10000;
	data_in <= 24'b010111100011111100010011;
#10000;
	data_in <= 24'b010111010011111000010001;
#10000;
	data_in <= 24'b010111000011110100010000;
#10000;
	data_in <= 24'b010110110011110100001111;
#10000;
	data_in <= 24'b010110100011101100001110;
#10000;
	data_in <= 24'b010110100011101000001101;
#10000;
	data_in <= 24'b010110000011100000001011;
#10000;
	data_in <= 24'b011000010100001100010110;
#10000;
	data_in <= 24'b011000000100001000010101;
#10000;
	data_in <= 24'b010111110100000000010100;
#10000;
	data_in <= 24'b010111100011111100010010;
#10000;
	data_in <= 24'b010111010011111000010001;
#10000;
	data_in <= 24'b010110110011110100010000;
#10000;
	data_in <= 24'b010110100011101100001111;
#10000;
	data_in <= 24'b010110100011101000001110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010110110011101100001111;
#10000;
	data_in <= 24'b010111000011110100010000;
#10000;
	data_in <= 24'b010111010011111000010010;
#10000;
	data_in <= 24'b010111110011111100010100;
#10000;
	data_in <= 24'b011000000100000000010101;
#10000;
	data_in <= 24'b011000010100001000010110;
#10000;
	data_in <= 24'b011000010100001100010110;
#10000;
	data_in <= 24'b011000100100010000011001;
#10000;
	data_in <= 24'b010111000011110100010000;
#10000;
	data_in <= 24'b010111100011111100010010;
#10000;
	data_in <= 24'b011000010100000000010011;
#10000;
	data_in <= 24'b011000010100000000010101;
#10000;
	data_in <= 24'b011000110100001000010111;
#10000;
	data_in <= 24'b011000110100001100010111;
#10000;
	data_in <= 24'b011001000100010000011001;
#10000;
	data_in <= 24'b011001010100011000011010;
#10000;
	data_in <= 24'b010111110100000000010011;
#10000;
	data_in <= 24'b011000010100000000010011;
#10000;
	data_in <= 24'b011000110100001000010110;
#10000;
	data_in <= 24'b011000110100001000010111;
#10000;
	data_in <= 24'b011001000100010000011000;
#10000;
	data_in <= 24'b011001010100010100011010;
#10000;
	data_in <= 24'b011001100100011000011011;
#10000;
	data_in <= 24'b011001110100011100011100;
#10000;
	data_in <= 24'b011000000100001000010101;
#10000;
	data_in <= 24'b011000100100001100010110;
#10000;
	data_in <= 24'b011001000100010000011000;
#10000;
	data_in <= 24'b011001010100010100011010;
#10000;
	data_in <= 24'b011001100100011000011011;
#10000;
	data_in <= 24'b011001110100100000011101;
#10000;
	data_in <= 24'b011010000100100100011110;
#10000;
	data_in <= 24'b011010010100101000100000;
#10000;
	data_in <= 24'b011000100100001100010110;
#10000;
	data_in <= 24'b011000110100010000011000;
#10000;
	data_in <= 24'b011001000100010100011001;
#10000;
	data_in <= 24'b011001010100011100011011;
#10000;
	data_in <= 24'b011001110100100100011101;
#10000;
	data_in <= 24'b011010010100101000011111;
#10000;
	data_in <= 24'b011010100100101100100001;
#10000;
	data_in <= 24'b011010110100110000100010;
#10000;
	data_in <= 24'b011001000100010100011000;
#10000;
	data_in <= 24'b011001010100011000011010;
#10000;
	data_in <= 24'b011001100100011100011011;
#10000;
	data_in <= 24'b011010000100100100011101;
#10000;
	data_in <= 24'b011010010100101100011111;
#10000;
	data_in <= 24'b011010100100110000100000;
#10000;
	data_in <= 24'b011011000100110100100011;
#10000;
	data_in <= 24'b011011010100111100100100;
#10000;
	data_in <= 24'b011001010100011000011010;
#10000;
	data_in <= 24'b011001110100100000011100;
#10000;
	data_in <= 24'b011010010100100100011110;
#10000;
	data_in <= 24'b011010100100110000100000;
#10000;
	data_in <= 24'b011010110100110100100001;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011011010101000000100101;
#10000;
	data_in <= 24'b011011110101000100100110;
#10000;
	data_in <= 24'b011001110100011100011100;
#10000;
	data_in <= 24'b011010010100100100011110;
#10000;
	data_in <= 24'b011010100100101100100001;
#10000;
	data_in <= 24'b011010110100110100100010;
#10000;
	data_in <= 24'b011011010100111100100100;
#10000;
	data_in <= 24'b011011100101000000100110;
#10000;
	data_in <= 24'b011011110101001000100111;
#10000;
	data_in <= 24'b011100010101010000101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000110100010100011010;
#10000;
	data_in <= 24'b011001000100011000011011;
#10000;
	data_in <= 24'b011001000100011000011100;
#10000;
	data_in <= 24'b011001010100011100011110;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001100100101000100000;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011010000100101100100010;
#10000;
	data_in <= 24'b011001010100011000011100;
#10000;
	data_in <= 24'b011001100100011100011101;
#10000;
	data_in <= 24'b011001110100100000011110;
#10000;
	data_in <= 24'b011010000100101000011111;
#10000;
	data_in <= 24'b011010000100101000100001;
#10000;
	data_in <= 24'b011010100100101100100010;
#10000;
	data_in <= 24'b011011000100110100100011;
#10000;
	data_in <= 24'b011011000100111000100100;
#10000;
	data_in <= 24'b011010000100100100011111;
#10000;
	data_in <= 24'b011010010100101100100000;
#10000;
	data_in <= 24'b011010010100110000100000;
#10000;
	data_in <= 24'b011010100100110000100010;
#10000;
	data_in <= 24'b011010110100110100100011;
#10000;
	data_in <= 24'b011011010100111000100100;
#10000;
	data_in <= 24'b011011010100111100100101;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011010100100110000100010;
#10000;
	data_in <= 24'b011010110100111000100011;
#10000;
	data_in <= 24'b011011000100111100100100;
#10000;
	data_in <= 24'b011011000100111100100101;
#10000;
	data_in <= 24'b011011100101000000100111;
#10000;
	data_in <= 24'b011011110101001000101000;
#10000;
	data_in <= 24'b011011110101001100101001;
#10000;
	data_in <= 24'b011100000101010000101010;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011011010100111100100101;
#10000;
	data_in <= 24'b011011100101000100100111;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011100000101001100101001;
#10000;
	data_in <= 24'b011100010101010000101011;
#10000;
	data_in <= 24'b011100100101010100101100;
#10000;
	data_in <= 24'b011100110101011100101100;
#10000;
	data_in <= 24'b011011100101000000100110;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011100010101001100101001;
#10000;
	data_in <= 24'b011100100101010100101011;
#10000;
	data_in <= 24'b011100110101011000101100;
#10000;
	data_in <= 24'b011101000101011100101101;
#10000;
	data_in <= 24'b011101010101100000101111;
#10000;
	data_in <= 24'b011101010101100100110000;
#10000;
	data_in <= 24'b011100000101001100101001;
#10000;
	data_in <= 24'b011100110101010000101011;
#10000;
	data_in <= 24'b011101000101011000101100;
#10000;
	data_in <= 24'b011101000101100000101110;
#10000;
	data_in <= 24'b011101100101100100101111;
#10000;
	data_in <= 24'b011101100101100100110000;
#10000;
	data_in <= 24'b011101110101101000110010;
#10000;
	data_in <= 24'b011110000101101100110100;
#10000;
	data_in <= 24'b011101000101010100101100;
#10000;
	data_in <= 24'b011101010101011100101101;
#10000;
	data_in <= 24'b011101100101100100101110;
#10000;
	data_in <= 24'b011101110101101000110001;
#10000;
	data_in <= 24'b011110000101101100110010;
#10000;
	data_in <= 24'b011110010101110000110011;
#10000;
	data_in <= 24'b011110100101110100110101;
#10000;
	data_in <= 24'b011110110101111000110111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011010100100110000100011;
#10000;
	data_in <= 24'b011010100100110100100100;
#10000;
	data_in <= 24'b011010110100111000100101;
#10000;
	data_in <= 24'b011010110100111100100111;
#10000;
	data_in <= 24'b011011000101000000100111;
#10000;
	data_in <= 24'b011011000101000000100111;
#10000;
	data_in <= 24'b011011000101000000101000;
#10000;
	data_in <= 24'b011011010101000100101001;
#10000;
	data_in <= 24'b011011010100111100100101;
#10000;
	data_in <= 24'b011011010100111100100111;
#10000;
	data_in <= 24'b011011100101000000100111;
#10000;
	data_in <= 24'b011011100101000100101000;
#10000;
	data_in <= 24'b011011110101001000101001;
#10000;
	data_in <= 24'b011011110101001100101010;
#10000;
	data_in <= 24'b011011110101001100101010;
#10000;
	data_in <= 24'b011100000101010000101011;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011100000101001000101001;
#10000;
	data_in <= 24'b011100000101001000101010;
#10000;
	data_in <= 24'b011100010101001100101011;
#10000;
	data_in <= 24'b011100010101010000101100;
#10000;
	data_in <= 24'b011100100101011000101101;
#10000;
	data_in <= 24'b011100100101011100101110;
#10000;
	data_in <= 24'b011100110101011000101111;
#10000;
	data_in <= 24'b011100100101010100101011;
#10000;
	data_in <= 24'b011100100101010100101011;
#10000;
	data_in <= 24'b011100110101011000101101;
#10000;
	data_in <= 24'b011101000101011100101111;
#10000;
	data_in <= 24'b011101010101100000101111;
#10000;
	data_in <= 24'b011101010101100100110000;
#10000;
	data_in <= 24'b011101010101101000110001;
#10000;
	data_in <= 24'b011101100101101100110010;
#10000;
	data_in <= 24'b011101010101100000101110;
#10000;
	data_in <= 24'b011101010101100000101111;
#10000;
	data_in <= 24'b011101100101100100110000;
#10000;
	data_in <= 24'b011101100101101000110001;
#10000;
	data_in <= 24'b011101110101101100110010;
#10000;
	data_in <= 24'b011101110101110000110011;
#10000;
	data_in <= 24'b011110000101110100110101;
#10000;
	data_in <= 24'b011110000101110100110101;
#10000;
	data_in <= 24'b011101100101101000110001;
#10000;
	data_in <= 24'b011110000101101100110010;
#10000;
	data_in <= 24'b011110000101110000110010;
#10000;
	data_in <= 24'b011110010101110100110100;
#10000;
	data_in <= 24'b011110100101111000110101;
#10000;
	data_in <= 24'b011110100101111000110110;
#10000;
	data_in <= 24'b011110110101111100110111;
#10000;
	data_in <= 24'b011110110110000000111000;
#10000;
	data_in <= 24'b011110010101110100110100;
#10000;
	data_in <= 24'b011110100101111000110101;
#10000;
	data_in <= 24'b011110110101111100110111;
#10000;
	data_in <= 24'b011111000110000000111001;
#10000;
	data_in <= 24'b011111010110000100111010;
#10000;
	data_in <= 24'b011111100110000100111010;
#10000;
	data_in <= 24'b011111110110001100111011;
#10000;
	data_in <= 24'b011111110110010000111101;
#10000;
	data_in <= 24'b011111000110000000111000;
#10000;
	data_in <= 24'b011111000110001000111001;
#10000;
	data_in <= 24'b011111110110001100111100;
#10000;
	data_in <= 24'b011111110110010000111100;
#10000;
	data_in <= 24'b011111110110010000111101;
#10000;
	data_in <= 24'b100000100110010100111111;
#10000;
	data_in <= 24'b100000100110011000111111;
#10000;
	data_in <= 24'b100000100110011101000000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011010101000100101001;
#10000;
	data_in <= 24'b011011010101001000101001;
#10000;
	data_in <= 24'b011011010101001000101011;
#10000;
	data_in <= 24'b011011110101010000101011;
#10000;
	data_in <= 24'b011011110101010000101100;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011100000101010000101100;
#10000;
	data_in <= 24'b011100000101010000101101;
#10000;
	data_in <= 24'b011100010101010100101110;
#10000;
	data_in <= 24'b011100100101010100101110;
#10000;
	data_in <= 24'b011100100101011000101110;
#10000;
	data_in <= 24'b011100100101011000101110;
#10000;
	data_in <= 24'b011100110101011000101111;
#10000;
	data_in <= 24'b011100100101011100101111;
#10000;
	data_in <= 24'b011100110101011100110000;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011101010101100100110001;
#10000;
	data_in <= 24'b011101010101100100110001;
#10000;
	data_in <= 24'b011101100101101000110011;
#10000;
	data_in <= 24'b011101110101101100110100;
#10000;
	data_in <= 24'b011101100101101100110011;
#10000;
	data_in <= 24'b011101100101101100110100;
#10000;
	data_in <= 24'b011101110101101100110100;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011110000101110100110110;
#10000;
	data_in <= 24'b011110010101111000110110;
#10000;
	data_in <= 24'b011110100101111100110111;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110000101110100110101;
#10000;
	data_in <= 24'b011110010101111000110110;
#10000;
	data_in <= 24'b011110100101111100111000;
#10000;
	data_in <= 24'b011110110101111100111001;
#10000;
	data_in <= 24'b011111000110000000111001;
#10000;
	data_in <= 24'b011111000110000100111001;
#10000;
	data_in <= 24'b011111000110000100111001;
#10000;
	data_in <= 24'b011111000110000100111010;
#10000;
	data_in <= 24'b011111000110000100111001;
#10000;
	data_in <= 24'b011111010110001000111010;
#10000;
	data_in <= 24'b011111100110001100111011;
#10000;
	data_in <= 24'b011111100110001100111100;
#10000;
	data_in <= 24'b011111110110001100111100;
#10000;
	data_in <= 24'b011111110110010000111100;
#10000;
	data_in <= 24'b011111110110010100111101;
#10000;
	data_in <= 24'b100000000110010100111110;
#10000;
	data_in <= 24'b100000000110010100111101;
#10000;
	data_in <= 24'b100000010110011000111110;
#10000;
	data_in <= 24'b100000010110011000111111;
#10000;
	data_in <= 24'b100000010110011001000000;
#10000;
	data_in <= 24'b100000100110011001000001;
#10000;
	data_in <= 24'b100000110110011101000001;
#10000;
	data_in <= 24'b100000110110100001000001;
#10000;
	data_in <= 24'b100000110110100001000010;
#10000;
	data_in <= 24'b100000110110100001000001;
#10000;
	data_in <= 24'b100000110110100001000010;
#10000;
	data_in <= 24'b100000110110100101000011;
#10000;
	data_in <= 24'b100001000110100101000100;
#10000;
	data_in <= 24'b100001010110101001000101;
#10000;
	data_in <= 24'b100001100110101001000101;
#10000;
	data_in <= 24'b100001100110101101000110;
#10000;
	data_in <= 24'b100001110110110001000110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011100000101010000101110;
#10000;
	data_in <= 24'b011100000101010000101110;
#10000;
	data_in <= 24'b011100000101010100101110;
#10000;
	data_in <= 24'b011100000101010100101110;
#10000;
	data_in <= 24'b011100000101011000101111;
#10000;
	data_in <= 24'b011100010101011000101111;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011000101111;
#10000;
	data_in <= 24'b011100110101011000110000;
#10000;
	data_in <= 24'b011100110101011100110001;
#10000;
	data_in <= 24'b011101000101100000110010;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011101000101100100110010;
#10000;
	data_in <= 24'b011101000101100100110010;
#10000;
	data_in <= 24'b011101000101100100110010;
#10000;
	data_in <= 24'b011101110101101000110011;
#10000;
	data_in <= 24'b011101110101101100110100;
#10000;
	data_in <= 24'b011101110101101100110101;
#10000;
	data_in <= 24'b011101110101101100110101;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011110100101111000110111;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011111010110001000111011;
#10000;
	data_in <= 24'b011111010110001000111011;
#10000;
	data_in <= 24'b011111010110001000111100;
#10000;
	data_in <= 24'b011111010110001000111101;
#10000;
	data_in <= 24'b011111010110001000111101;
#10000;
	data_in <= 24'b011111010110001100111101;
#10000;
	data_in <= 24'b011111010110001100111101;
#10000;
	data_in <= 24'b011111010110001100111101;
#10000;
	data_in <= 24'b100000000110010100111111;
#10000;
	data_in <= 24'b100000000110010100111111;
#10000;
	data_in <= 24'b100000000110010100111111;
#10000;
	data_in <= 24'b100000000110010101000000;
#10000;
	data_in <= 24'b100000000110011001000000;
#10000;
	data_in <= 24'b100000000110011101000000;
#10000;
	data_in <= 24'b100000000110011001000000;
#10000;
	data_in <= 24'b100000000110011101000001;
#10000;
	data_in <= 24'b100000110110100001000010;
#10000;
	data_in <= 24'b100000110110100001000011;
#10000;
	data_in <= 24'b100000110110100101000100;
#10000;
	data_in <= 24'b100000110110101001000100;
#10000;
	data_in <= 24'b100000110110101001000100;
#10000;
	data_in <= 24'b100000110110101101000101;
#10000;
	data_in <= 24'b100000110110101101000101;
#10000;
	data_in <= 24'b100000110110101101000101;
#10000;
	data_in <= 24'b100001110110110001000111;
#10000;
	data_in <= 24'b100001110110110101001000;
#10000;
	data_in <= 24'b100001110110110001001000;
#10000;
	data_in <= 24'b100001110110110101001000;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
	data_in <= 24'b100001100110110101001000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011101010101100100110011;
#10000;
	data_in <= 24'b011101010101100100110010;
#10000;
	data_in <= 24'b011101010101100100110010;
#10000;
	data_in <= 24'b011101010101100100110010;
#10000;
	data_in <= 24'b011101010101100100110011;
#10000;
	data_in <= 24'b011101010101101000110100;
#10000;
	data_in <= 24'b011101010101101000110011;
#10000;
	data_in <= 24'b011101010101101000110011;
#10000;
	data_in <= 24'b011110000101110000110110;
#10000;
	data_in <= 24'b011110000101110000110111;
#10000;
	data_in <= 24'b011110000101110000110111;
#10000;
	data_in <= 24'b011110000101110000110110;
#10000;
	data_in <= 24'b011110000101110100110111;
#10000;
	data_in <= 24'b011110000101110100111000;
#10000;
	data_in <= 24'b011110000101110100111000;
#10000;
	data_in <= 24'b011110000101110100111000;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b100000010110011001000010;
#10000;
	data_in <= 24'b100000010110011101000010;
#10000;
	data_in <= 24'b100000010110011101000010;
#10000;
	data_in <= 24'b100000010110100001000010;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100001000110101101000101;
#10000;
	data_in <= 24'b100001000110101001000110;
#10000;
	data_in <= 24'b100001000110101101000101;
#10000;
	data_in <= 24'b100001000110110001000101;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
	data_in <= 24'b100010000110110101001010;
#10000;
	data_in <= 24'b100001110110111001001010;
#10000;
	data_in <= 24'b100010000110111001001001;
#10000;
	data_in <= 24'b100010000110111001001010;
#10000;
	data_in <= 24'b100010000110111001001011;
#10000;
	data_in <= 24'b100010000110111001001011;
#10000;
	data_in <= 24'b100010000110111001001011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011100100101011100110001;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011101010101101000110011;
#10000;
	data_in <= 24'b011101010101101000110011;
#10000;
	data_in <= 24'b011101010101101000110100;
#10000;
	data_in <= 24'b011101010101100100110011;
#10000;
	data_in <= 24'b011101010101100100110010;
#10000;
	data_in <= 24'b011101010101100100110010;
#10000;
	data_in <= 24'b011101010101100100110010;
#10000;
	data_in <= 24'b011101010101100100110011;
#10000;
	data_in <= 24'b011110000101110100111000;
#10000;
	data_in <= 24'b011110000101110100111000;
#10000;
	data_in <= 24'b011110000101110100111000;
#10000;
	data_in <= 24'b011110000101110100110111;
#10000;
	data_in <= 24'b011110000101110000110110;
#10000;
	data_in <= 24'b011110000101110000110111;
#10000;
	data_in <= 24'b011110000101110000110111;
#10000;
	data_in <= 24'b011110000101110000110110;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011110110110000000111011;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011110110101111100111010;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b011111100110010000111111;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b011111100110001100111110;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100000010110100001000011;
#10000;
	data_in <= 24'b100000010110100001000010;
#10000;
	data_in <= 24'b100000010110011101000010;
#10000;
	data_in <= 24'b100000010110011101000010;
#10000;
	data_in <= 24'b100000010110011001000010;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001000110101101000110;
#10000;
	data_in <= 24'b100001000110110001000101;
#10000;
	data_in <= 24'b100001000110101101000101;
#10000;
	data_in <= 24'b100001000110101001000110;
#10000;
	data_in <= 24'b100001000110101101000101;
#10000;
	data_in <= 24'b100010000110111001001011;
#10000;
	data_in <= 24'b100010000110111001001011;
#10000;
	data_in <= 24'b100010000110111001001011;
#10000;
	data_in <= 24'b100010000110111001001010;
#10000;
	data_in <= 24'b100010000110111001001001;
#10000;
	data_in <= 24'b100001110110111001001010;
#10000;
	data_in <= 24'b100010000110110101001010;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100100101011000110000;
#10000;
	data_in <= 24'b011100010101011000101111;
#10000;
	data_in <= 24'b011100000101011000101111;
#10000;
	data_in <= 24'b011100000101010100101110;
#10000;
	data_in <= 24'b011100000101010100101110;
#10000;
	data_in <= 24'b011100000101010000101110;
#10000;
	data_in <= 24'b011100000101010000101110;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011101000101100100110010;
#10000;
	data_in <= 24'b011101000101100100110010;
#10000;
	data_in <= 24'b011101000101100100110010;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011101000101100000110010;
#10000;
	data_in <= 24'b011100110101011100110001;
#10000;
	data_in <= 24'b011100110101011000110000;
#10000;
	data_in <= 24'b011100100101011000101111;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101101100110101;
#10000;
	data_in <= 24'b011101110101101100110101;
#10000;
	data_in <= 24'b011101110101101100110100;
#10000;
	data_in <= 24'b011101110101101000110011;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011110100101111100111001;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110100101111000110111;
#10000;
	data_in <= 24'b011111010110001100111101;
#10000;
	data_in <= 24'b011111010110001100111101;
#10000;
	data_in <= 24'b011111010110001100111101;
#10000;
	data_in <= 24'b011111010110001000111101;
#10000;
	data_in <= 24'b011111010110001000111101;
#10000;
	data_in <= 24'b011111010110001000111100;
#10000;
	data_in <= 24'b011111010110001000111011;
#10000;
	data_in <= 24'b011111010110001000111011;
#10000;
	data_in <= 24'b100000000110011101000001;
#10000;
	data_in <= 24'b100000000110011001000000;
#10000;
	data_in <= 24'b100000000110011101000000;
#10000;
	data_in <= 24'b100000000110011001000000;
#10000;
	data_in <= 24'b100000000110010101000000;
#10000;
	data_in <= 24'b100000000110010100111111;
#10000;
	data_in <= 24'b100000000110010100111111;
#10000;
	data_in <= 24'b100000000110010100111111;
#10000;
	data_in <= 24'b100000110110101101000101;
#10000;
	data_in <= 24'b100000110110101101000101;
#10000;
	data_in <= 24'b100000110110101101000101;
#10000;
	data_in <= 24'b100000110110101001000100;
#10000;
	data_in <= 24'b100000110110101001000100;
#10000;
	data_in <= 24'b100000110110100101000100;
#10000;
	data_in <= 24'b100000110110100001000011;
#10000;
	data_in <= 24'b100000110110100001000010;
#10000;
	data_in <= 24'b100001100110110101001000;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
	data_in <= 24'b100001110110110101001001;
#10000;
	data_in <= 24'b100001110110110101001000;
#10000;
	data_in <= 24'b100001110110110001001000;
#10000;
	data_in <= 24'b100001110110110101001000;
#10000;
	data_in <= 24'b100001110110110001000111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101101;
#10000;
	data_in <= 24'b011011110101010000101100;
#10000;
	data_in <= 24'b011011110101010000101011;
#10000;
	data_in <= 24'b011011010101001000101011;
#10000;
	data_in <= 24'b011011010101001000101001;
#10000;
	data_in <= 24'b011011010101000100101001;
#10000;
	data_in <= 24'b011100100101011100101111;
#10000;
	data_in <= 24'b011100110101011000101111;
#10000;
	data_in <= 24'b011100100101011000101110;
#10000;
	data_in <= 24'b011100100101011000101110;
#10000;
	data_in <= 24'b011100100101010100101110;
#10000;
	data_in <= 24'b011100010101010100101110;
#10000;
	data_in <= 24'b011100000101010000101101;
#10000;
	data_in <= 24'b011100000101010000101100;
#10000;
	data_in <= 24'b011101110101101100110100;
#10000;
	data_in <= 24'b011101100101101000110011;
#10000;
	data_in <= 24'b011101010101100100110001;
#10000;
	data_in <= 24'b011101010101100100110001;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011101000101100000110001;
#10000;
	data_in <= 24'b011100110101011100110000;
#10000;
	data_in <= 24'b011110100101111000111000;
#10000;
	data_in <= 24'b011110100101111100110111;
#10000;
	data_in <= 24'b011110010101111000110110;
#10000;
	data_in <= 24'b011110000101110100110110;
#10000;
	data_in <= 24'b011101110101110000110101;
#10000;
	data_in <= 24'b011101110101101100110100;
#10000;
	data_in <= 24'b011101100101101100110100;
#10000;
	data_in <= 24'b011101100101101100110011;
#10000;
	data_in <= 24'b011111000110000100111010;
#10000;
	data_in <= 24'b011111000110000100111001;
#10000;
	data_in <= 24'b011111000110000100111001;
#10000;
	data_in <= 24'b011111000110000000111001;
#10000;
	data_in <= 24'b011110110101111100111001;
#10000;
	data_in <= 24'b011110100101111100111000;
#10000;
	data_in <= 24'b011110010101111000110110;
#10000;
	data_in <= 24'b011110000101110100110101;
#10000;
	data_in <= 24'b100000000110010100111110;
#10000;
	data_in <= 24'b011111110110010100111101;
#10000;
	data_in <= 24'b011111110110010000111100;
#10000;
	data_in <= 24'b011111110110001100111100;
#10000;
	data_in <= 24'b011111100110001100111100;
#10000;
	data_in <= 24'b011111100110001100111011;
#10000;
	data_in <= 24'b011111010110001000111010;
#10000;
	data_in <= 24'b011111000110000100111001;
#10000;
	data_in <= 24'b100000110110100001000010;
#10000;
	data_in <= 24'b100000110110100001000001;
#10000;
	data_in <= 24'b100000110110011101000001;
#10000;
	data_in <= 24'b100000100110011001000001;
#10000;
	data_in <= 24'b100000010110011001000000;
#10000;
	data_in <= 24'b100000010110011000111111;
#10000;
	data_in <= 24'b100000010110011000111110;
#10000;
	data_in <= 24'b100000000110010100111101;
#10000;
	data_in <= 24'b100001110110110001000110;
#10000;
	data_in <= 24'b100001100110101101000110;
#10000;
	data_in <= 24'b100001100110101001000101;
#10000;
	data_in <= 24'b100001010110101001000101;
#10000;
	data_in <= 24'b100001000110100101000100;
#10000;
	data_in <= 24'b100000110110100101000011;
#10000;
	data_in <= 24'b100000110110100001000010;
#10000;
	data_in <= 24'b100000110110100001000001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011010101000100101001;
#10000;
	data_in <= 24'b011011000101000000101000;
#10000;
	data_in <= 24'b011011000101000000100111;
#10000;
	data_in <= 24'b011011000101000000100111;
#10000;
	data_in <= 24'b011010110100111100100111;
#10000;
	data_in <= 24'b011010110100111000100101;
#10000;
	data_in <= 24'b011010100100110100100100;
#10000;
	data_in <= 24'b011010100100110000100011;
#10000;
	data_in <= 24'b011100000101010000101011;
#10000;
	data_in <= 24'b011011110101001100101010;
#10000;
	data_in <= 24'b011011110101001100101010;
#10000;
	data_in <= 24'b011011110101001000101001;
#10000;
	data_in <= 24'b011011100101000100101000;
#10000;
	data_in <= 24'b011011100101000000100111;
#10000;
	data_in <= 24'b011011010100111100100111;
#10000;
	data_in <= 24'b011011010100111100100101;
#10000;
	data_in <= 24'b011100110101011000101111;
#10000;
	data_in <= 24'b011100100101011100101110;
#10000;
	data_in <= 24'b011100100101011000101101;
#10000;
	data_in <= 24'b011100010101010000101100;
#10000;
	data_in <= 24'b011100010101001100101011;
#10000;
	data_in <= 24'b011100000101001000101010;
#10000;
	data_in <= 24'b011100000101001000101001;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011101100101101100110010;
#10000;
	data_in <= 24'b011101010101101000110001;
#10000;
	data_in <= 24'b011101010101100100110000;
#10000;
	data_in <= 24'b011101010101100000101111;
#10000;
	data_in <= 24'b011101000101011100101111;
#10000;
	data_in <= 24'b011100110101011000101101;
#10000;
	data_in <= 24'b011100100101010100101011;
#10000;
	data_in <= 24'b011100100101010100101011;
#10000;
	data_in <= 24'b011110000101110100110101;
#10000;
	data_in <= 24'b011110000101110100110101;
#10000;
	data_in <= 24'b011101110101110000110011;
#10000;
	data_in <= 24'b011101110101101100110010;
#10000;
	data_in <= 24'b011101100101101000110001;
#10000;
	data_in <= 24'b011101100101100100110000;
#10000;
	data_in <= 24'b011101010101100000101111;
#10000;
	data_in <= 24'b011101010101100000101110;
#10000;
	data_in <= 24'b011110110110000000111000;
#10000;
	data_in <= 24'b011110110101111100110111;
#10000;
	data_in <= 24'b011110100101111000110110;
#10000;
	data_in <= 24'b011110100101111000110101;
#10000;
	data_in <= 24'b011110010101110100110100;
#10000;
	data_in <= 24'b011110000101110000110010;
#10000;
	data_in <= 24'b011110000101101100110010;
#10000;
	data_in <= 24'b011101100101101000110001;
#10000;
	data_in <= 24'b011111110110010000111101;
#10000;
	data_in <= 24'b011111110110001100111011;
#10000;
	data_in <= 24'b011111100110000100111010;
#10000;
	data_in <= 24'b011111010110000100111010;
#10000;
	data_in <= 24'b011111000110000000111001;
#10000;
	data_in <= 24'b011110110101111100110111;
#10000;
	data_in <= 24'b011110100101111000110101;
#10000;
	data_in <= 24'b011110010101110100110100;
#10000;
	data_in <= 24'b100000100110011101000000;
#10000;
	data_in <= 24'b100000100110011000111111;
#10000;
	data_in <= 24'b100000100110010100111111;
#10000;
	data_in <= 24'b011111110110010000111101;
#10000;
	data_in <= 24'b011111110110010000111100;
#10000;
	data_in <= 24'b011111110110001100111100;
#10000;
	data_in <= 24'b011111000110001000111001;
#10000;
	data_in <= 24'b011111000110000000111000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011010000100101100100010;
#10000;
	data_in <= 24'b011001110100101100100001;
#10000;
	data_in <= 24'b011001100100101000100000;
#10000;
	data_in <= 24'b011001010100100000011110;
#10000;
	data_in <= 24'b011001010100011100011110;
#10000;
	data_in <= 24'b011001000100011000011100;
#10000;
	data_in <= 24'b011001000100011000011011;
#10000;
	data_in <= 24'b011000110100010100011010;
#10000;
	data_in <= 24'b011011000100111000100100;
#10000;
	data_in <= 24'b011011000100110100100011;
#10000;
	data_in <= 24'b011010100100101100100010;
#10000;
	data_in <= 24'b011010000100101000100001;
#10000;
	data_in <= 24'b011010000100101000011111;
#10000;
	data_in <= 24'b011001110100100000011110;
#10000;
	data_in <= 24'b011001100100011100011101;
#10000;
	data_in <= 24'b011001010100011000011100;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011011010100111100100101;
#10000;
	data_in <= 24'b011011010100111000100100;
#10000;
	data_in <= 24'b011010110100110100100011;
#10000;
	data_in <= 24'b011010100100110000100010;
#10000;
	data_in <= 24'b011010010100110000100000;
#10000;
	data_in <= 24'b011010010100101100100000;
#10000;
	data_in <= 24'b011010000100100100011111;
#10000;
	data_in <= 24'b011100000101010000101010;
#10000;
	data_in <= 24'b011011110101001100101001;
#10000;
	data_in <= 24'b011011110101001000101000;
#10000;
	data_in <= 24'b011011100101000000100111;
#10000;
	data_in <= 24'b011011000100111100100101;
#10000;
	data_in <= 24'b011011000100111100100100;
#10000;
	data_in <= 24'b011010110100111000100011;
#10000;
	data_in <= 24'b011010100100110000100010;
#10000;
	data_in <= 24'b011100110101011100101100;
#10000;
	data_in <= 24'b011100100101010100101100;
#10000;
	data_in <= 24'b011100010101010000101011;
#10000;
	data_in <= 24'b011100000101001100101001;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011011100101000100100111;
#10000;
	data_in <= 24'b011011010100111100100101;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011101010101100100110000;
#10000;
	data_in <= 24'b011101010101100000101111;
#10000;
	data_in <= 24'b011101000101011100101101;
#10000;
	data_in <= 24'b011100110101011000101100;
#10000;
	data_in <= 24'b011100100101010100101011;
#10000;
	data_in <= 24'b011100010101001100101001;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011011100101000000100110;
#10000;
	data_in <= 24'b011110000101101100110100;
#10000;
	data_in <= 24'b011101110101101000110010;
#10000;
	data_in <= 24'b011101100101100100110000;
#10000;
	data_in <= 24'b011101100101100100101111;
#10000;
	data_in <= 24'b011101000101100000101110;
#10000;
	data_in <= 24'b011101000101011000101100;
#10000;
	data_in <= 24'b011100110101010000101011;
#10000;
	data_in <= 24'b011100000101001100101001;
#10000;
	data_in <= 24'b011110110101111000110111;
#10000;
	data_in <= 24'b011110100101110100110101;
#10000;
	data_in <= 24'b011110010101110000110011;
#10000;
	data_in <= 24'b011110000101101100110010;
#10000;
	data_in <= 24'b011101110101101000110001;
#10000;
	data_in <= 24'b011101100101100100101110;
#10000;
	data_in <= 24'b011101010101011100101101;
#10000;
	data_in <= 24'b011101000101010100101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000100100010000011001;
#10000;
	data_in <= 24'b011000010100001100010110;
#10000;
	data_in <= 24'b011000010100001000010110;
#10000;
	data_in <= 24'b011000000100000000010101;
#10000;
	data_in <= 24'b010111110011111100010100;
#10000;
	data_in <= 24'b010111010011111000010010;
#10000;
	data_in <= 24'b010111000011110100010000;
#10000;
	data_in <= 24'b010110110011101100001111;
#10000;
	data_in <= 24'b011001010100011000011010;
#10000;
	data_in <= 24'b011001000100010000011001;
#10000;
	data_in <= 24'b011000110100001100010111;
#10000;
	data_in <= 24'b011000110100001000010111;
#10000;
	data_in <= 24'b011000010100000000010101;
#10000;
	data_in <= 24'b011000010100000000010011;
#10000;
	data_in <= 24'b010111100011111100010010;
#10000;
	data_in <= 24'b010111000011110100010000;
#10000;
	data_in <= 24'b011001110100011100011100;
#10000;
	data_in <= 24'b011001100100011000011011;
#10000;
	data_in <= 24'b011001010100010100011010;
#10000;
	data_in <= 24'b011001000100010000011000;
#10000;
	data_in <= 24'b011000110100001000010111;
#10000;
	data_in <= 24'b011000110100001000010110;
#10000;
	data_in <= 24'b011000010100000000010011;
#10000;
	data_in <= 24'b010111110100000000010011;
#10000;
	data_in <= 24'b011010010100101000100000;
#10000;
	data_in <= 24'b011010000100100100011110;
#10000;
	data_in <= 24'b011001110100100000011101;
#10000;
	data_in <= 24'b011001100100011000011011;
#10000;
	data_in <= 24'b011001010100010100011010;
#10000;
	data_in <= 24'b011001000100010000011000;
#10000;
	data_in <= 24'b011000100100001100010110;
#10000;
	data_in <= 24'b011000000100001000010101;
#10000;
	data_in <= 24'b011010110100110000100010;
#10000;
	data_in <= 24'b011010100100101100100001;
#10000;
	data_in <= 24'b011010010100101000011111;
#10000;
	data_in <= 24'b011001110100100100011101;
#10000;
	data_in <= 24'b011001010100011100011011;
#10000;
	data_in <= 24'b011001000100010100011001;
#10000;
	data_in <= 24'b011000110100010000011000;
#10000;
	data_in <= 24'b011000100100001100010110;
#10000;
	data_in <= 24'b011011010100111100100100;
#10000;
	data_in <= 24'b011011000100110100100011;
#10000;
	data_in <= 24'b011010100100110000100000;
#10000;
	data_in <= 24'b011010010100101100011111;
#10000;
	data_in <= 24'b011010000100100100011101;
#10000;
	data_in <= 24'b011001100100011100011011;
#10000;
	data_in <= 24'b011001010100011000011010;
#10000;
	data_in <= 24'b011001000100010100011000;
#10000;
	data_in <= 24'b011011110101000100100110;
#10000;
	data_in <= 24'b011011010101000000100101;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011010110100110100100001;
#10000;
	data_in <= 24'b011010100100110000100000;
#10000;
	data_in <= 24'b011010010100100100011110;
#10000;
	data_in <= 24'b011001110100100000011100;
#10000;
	data_in <= 24'b011001010100011000011010;
#10000;
	data_in <= 24'b011100010101010000101001;
#10000;
	data_in <= 24'b011011110101001000100111;
#10000;
	data_in <= 24'b011011100101000000100110;
#10000;
	data_in <= 24'b011011010100111100100100;
#10000;
	data_in <= 24'b011010110100110100100010;
#10000;
	data_in <= 24'b011010100100101100100001;
#10000;
	data_in <= 24'b011010010100100100011110;
#10000;
	data_in <= 24'b011001110100011100011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011010010100101000011110;
#10000;
	data_in <= 24'b011010100100110000100000;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011011010100111100100100;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011100010101010000101001;
#10000;
	data_in <= 24'b011100100101011000101010;
#10000;
	data_in <= 24'b011101000101011100101100;
#10000;
	data_in <= 24'b011010110100110000100000;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011011100101000000100101;
#10000;
	data_in <= 24'b011100000101001000100111;
#10000;
	data_in <= 24'b011100010101010000101010;
#10000;
	data_in <= 24'b011100110101011100101011;
#10000;
	data_in <= 24'b011101000101100000101101;
#10000;
	data_in <= 24'b011101100101100100110000;
#10000;
	data_in <= 24'b011011010100111000100011;
#10000;
	data_in <= 24'b011011110101000000100101;
#10000;
	data_in <= 24'b011100000101001000100111;
#10000;
	data_in <= 24'b011100100101010000101001;
#10000;
	data_in <= 24'b011101000101011100101100;
#10000;
	data_in <= 24'b011101010101100100101110;
#10000;
	data_in <= 24'b011101110101101000110000;
#10000;
	data_in <= 24'b011110010101110000110010;
#10000;
	data_in <= 24'b011011110101000000100101;
#10000;
	data_in <= 24'b011100000101001100100111;
#10000;
	data_in <= 24'b011100100101010000101001;
#10000;
	data_in <= 24'b011101000101011000101011;
#10000;
	data_in <= 24'b011101100101100100101110;
#10000;
	data_in <= 24'b011110000101101100110001;
#10000;
	data_in <= 24'b011110100101110100110011;
#10000;
	data_in <= 24'b011111000101111100110101;
#10000;
	data_in <= 24'b011100010101001100101000;
#10000;
	data_in <= 24'b011100110101010100101010;
#10000;
	data_in <= 24'b011101010101011100101100;
#10000;
	data_in <= 24'b011101100101100100101111;
#10000;
	data_in <= 24'b011110000101101100110000;
#10000;
	data_in <= 24'b011110110101110100110011;
#10000;
	data_in <= 24'b011111010110000000110111;
#10000;
	data_in <= 24'b011111100110001000111000;
#10000;
	data_in <= 24'b011100110101010100101010;
#10000;
	data_in <= 24'b011101010101011100101100;
#10000;
	data_in <= 24'b011101110101100100101111;
#10000;
	data_in <= 24'b011110100101110000110010;
#10000;
	data_in <= 24'b011111000101111000110100;
#10000;
	data_in <= 24'b011111010110000000110110;
#10000;
	data_in <= 24'b100000000110001000111001;
#10000;
	data_in <= 24'b100000100110010100111011;
#10000;
	data_in <= 24'b011101010101011100101011;
#10000;
	data_in <= 24'b011101110101100100101101;
#10000;
	data_in <= 24'b011110100101110000110000;
#10000;
	data_in <= 24'b011111000101111100110100;
#10000;
	data_in <= 24'b011111010110000100110110;
#10000;
	data_in <= 24'b100000000110001000111001;
#10000;
	data_in <= 24'b100000100110010100111010;
#10000;
	data_in <= 24'b100001010110100000111110;
#10000;
	data_in <= 24'b011101110101100100101110;
#10000;
	data_in <= 24'b011110010101101100110001;
#10000;
	data_in <= 24'b011111000101111000110100;
#10000;
	data_in <= 24'b011111100110000000110111;
#10000;
	data_in <= 24'b100000000110001100111010;
#10000;
	data_in <= 24'b100000100110010000111011;
#10000;
	data_in <= 24'b100001010110011100111110;
#10000;
	data_in <= 24'b100001110110101001000010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011101100101100000101111;
#10000;
	data_in <= 24'b011101110101100100101111;
#10000;
	data_in <= 24'b011110000101110000110001;
#10000;
	data_in <= 24'b011110100101111000110011;
#10000;
	data_in <= 24'b011110110101111100110101;
#10000;
	data_in <= 24'b011111000110000000110111;
#10000;
	data_in <= 24'b011111010110000100111000;
#10000;
	data_in <= 24'b011111100110001100111001;
#10000;
	data_in <= 24'b011110000101101100110010;
#10000;
	data_in <= 24'b011110100101110100110011;
#10000;
	data_in <= 24'b011111000101111000110101;
#10000;
	data_in <= 24'b011111010110000000110110;
#10000;
	data_in <= 24'b011111100110001000111001;
#10000;
	data_in <= 24'b011111110110001100111011;
#10000;
	data_in <= 24'b100000000110010100111011;
#10000;
	data_in <= 24'b100000010110011000111101;
#10000;
	data_in <= 24'b011110100101111000110100;
#10000;
	data_in <= 24'b011111000110000000110111;
#10000;
	data_in <= 24'b011111100110001000111001;
#10000;
	data_in <= 24'b100000000110001100111010;
#10000;
	data_in <= 24'b100000000110010000111100;
#10000;
	data_in <= 24'b100000100110011000111110;
#10000;
	data_in <= 24'b100000110110100000111111;
#10000;
	data_in <= 24'b100001010110100101000001;
#10000;
	data_in <= 24'b011111100110000100110111;
#10000;
	data_in <= 24'b011111110110001100111010;
#10000;
	data_in <= 24'b100000010110010100111011;
#10000;
	data_in <= 24'b100000110110010100111101;
#10000;
	data_in <= 24'b100001000110100000111111;
#10000;
	data_in <= 24'b100001010110101001000001;
#10000;
	data_in <= 24'b100001100110101101000011;
#10000;
	data_in <= 24'b100001110110110001000100;
#10000;
	data_in <= 24'b100000000110010000111010;
#10000;
	data_in <= 24'b100000100110011000111101;
#10000;
	data_in <= 24'b100001000110011100111111;
#10000;
	data_in <= 24'b100001100110100101000001;
#10000;
	data_in <= 24'b100001110110101101000011;
#10000;
	data_in <= 24'b100010000110110101000101;
#10000;
	data_in <= 24'b100010100110111101000111;
#10000;
	data_in <= 24'b100010110111000001001000;
#10000;
	data_in <= 24'b100000110110011100111101;
#10000;
	data_in <= 24'b100001100110100101000000;
#10000;
	data_in <= 24'b100010000110101101000011;
#10000;
	data_in <= 24'b100010010110110001000100;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100011000111000101001000;
#10000;
	data_in <= 24'b100011010111001001001010;
#10000;
	data_in <= 24'b100011100111001101001100;
#10000;
	data_in <= 24'b100001100110101001000000;
#10000;
	data_in <= 24'b100010000110110001000010;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100011000110111101000111;
#10000;
	data_in <= 24'b100011010111001001001000;
#10000;
	data_in <= 24'b100011110111010001001011;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b100100100111011101001111;
#10000;
	data_in <= 24'b100010000110110001000011;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100011000111000001001001;
#10000;
	data_in <= 24'b100011100111001001001010;
#10000;
	data_in <= 24'b100100000111010101001101;
#10000;
	data_in <= 24'b100100100111011101001111;
#10000;
	data_in <= 24'b100101000111100001010000;
#10000;
	data_in <= 24'b100101010111101001010011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011111110110010000111011;
#10000;
	data_in <= 24'b011111110110010100111101;
#10000;
	data_in <= 24'b100000010110011100111110;
#10000;
	data_in <= 24'b100000100110011100111111;
#10000;
	data_in <= 24'b100001000110100001000000;
#10000;
	data_in <= 24'b100001010110100001000010;
#10000;
	data_in <= 24'b100001010110101001000010;
#10000;
	data_in <= 24'b100001100110110001000011;
#10000;
	data_in <= 24'b100000100110011100111111;
#10000;
	data_in <= 24'b100000110110100101000000;
#10000;
	data_in <= 24'b100001000110101001000010;
#10000;
	data_in <= 24'b100001110110101101000100;
#10000;
	data_in <= 24'b100010000110110001000101;
#10000;
	data_in <= 24'b100010000110110101000101;
#10000;
	data_in <= 24'b100010010110111001000110;
#10000;
	data_in <= 24'b100010010110111101001000;
#10000;
	data_in <= 24'b100001010110101001000010;
#10000;
	data_in <= 24'b100001100110101101000100;
#10000;
	data_in <= 24'b100010000110110101000110;
#10000;
	data_in <= 24'b100010100110111001001000;
#10000;
	data_in <= 24'b100010110110111101001001;
#10000;
	data_in <= 24'b100010110111000001001001;
#10000;
	data_in <= 24'b100011000111000101001010;
#10000;
	data_in <= 24'b100011010111001001001100;
#10000;
	data_in <= 24'b100010010110111001000110;
#10000;
	data_in <= 24'b100010100110111001001000;
#10000;
	data_in <= 24'b100011000111000001001001;
#10000;
	data_in <= 24'b100011000111001001001010;
#10000;
	data_in <= 24'b100011100111001101001100;
#10000;
	data_in <= 24'b100011110111010001001101;
#10000;
	data_in <= 24'b100100000111010101001110;
#10000;
	data_in <= 24'b100100000111011001010000;
#10000;
	data_in <= 24'b100011010111000101001010;
#10000;
	data_in <= 24'b100011100111001001001100;
#10000;
	data_in <= 24'b100011110111010101001110;
#10000;
	data_in <= 24'b100100000111011001001110;
#10000;
	data_in <= 24'b100100100111011101010000;
#10000;
	data_in <= 24'b100100110111100001010010;
#10000;
	data_in <= 24'b100100110111100001010011;
#10000;
	data_in <= 24'b100101000111101001010100;
#10000;
	data_in <= 24'b100100000111010101001110;
#10000;
	data_in <= 24'b100100010111011101010000;
#10000;
	data_in <= 24'b100100100111100101010001;
#10000;
	data_in <= 24'b100101000111101001010010;
#10000;
	data_in <= 24'b100101100111101101010100;
#10000;
	data_in <= 24'b100101110111110001010110;
#10000;
	data_in <= 24'b100101110111110001010110;
#10000;
	data_in <= 24'b100110000111110101010111;
#10000;
	data_in <= 24'b100100100111100101010001;
#10000;
	data_in <= 24'b100101000111101001010011;
#10000;
	data_in <= 24'b100101100111101101010100;
#10000;
	data_in <= 24'b100110000111110101010110;
#10000;
	data_in <= 24'b100110010111111001010111;
#10000;
	data_in <= 24'b100110100111111101011001;
#10000;
	data_in <= 24'b100110111000000001011010;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100101100111110001010101;
#10000;
	data_in <= 24'b100110000111110101010111;
#10000;
	data_in <= 24'b100110100111111101011001;
#10000;
	data_in <= 24'b100110101000000001011010;
#10000;
	data_in <= 24'b100111001000001001011100;
#10000;
	data_in <= 24'b100111101000001101011101;
#10000;
	data_in <= 24'b100111101000010001011110;
#10000;
	data_in <= 24'b100111111000010101011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100001100110110001000101;
#10000;
	data_in <= 24'b100001110110110101000110;
#10000;
	data_in <= 24'b100010000110111001000110;
#10000;
	data_in <= 24'b100010000110111001000111;
#10000;
	data_in <= 24'b100010010110111101001001;
#10000;
	data_in <= 24'b100010100111000001001001;
#10000;
	data_in <= 24'b100010100111000001001011;
#10000;
	data_in <= 24'b100010100111000101001011;
#10000;
	data_in <= 24'b100010100111000001001001;
#10000;
	data_in <= 24'b100010110111000101001010;
#10000;
	data_in <= 24'b100010110111000101001010;
#10000;
	data_in <= 24'b100010110111001001001011;
#10000;
	data_in <= 24'b100010110111001101001101;
#10000;
	data_in <= 24'b100011000111010001001101;
#10000;
	data_in <= 24'b100011010111010001001110;
#10000;
	data_in <= 24'b100011010111010101001110;
#10000;
	data_in <= 24'b100011010111001101001101;
#10000;
	data_in <= 24'b100011100111010001001110;
#10000;
	data_in <= 24'b100011100111010101001111;
#10000;
	data_in <= 24'b100011110111011001001111;
#10000;
	data_in <= 24'b100100000111011101010001;
#10000;
	data_in <= 24'b100100000111011101010010;
#10000;
	data_in <= 24'b100100010111100001010010;
#10000;
	data_in <= 24'b100100010111100001010011;
#10000;
	data_in <= 24'b100100010111100001010001;
#10000;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b100100110111101001010100;
#10000;
	data_in <= 24'b100100110111101001010100;
#10000;
	data_in <= 24'b100101000111101101010101;
#10000;
	data_in <= 24'b100101000111101101010101;
#10000;
	data_in <= 24'b100101010111110001010111;
#10000;
	data_in <= 24'b100101010111101101010101;
#10000;
	data_in <= 24'b100101010111110001010110;
#10000;
	data_in <= 24'b100101100111110101010111;
#10000;
	data_in <= 24'b100101100111110101011000;
#10000;
	data_in <= 24'b100101100111110101011001;
#10000;
	data_in <= 24'b100101110111111001011010;
#10000;
	data_in <= 24'b100110011000000001011011;
#10000;
	data_in <= 24'b100110011000000001011100;
#10000;
	data_in <= 24'b100110011000000001011010;
#10000;
	data_in <= 24'b100110101000000101011011;
#10000;
	data_in <= 24'b100110101000000101011100;
#10000;
	data_in <= 24'b100110111000001001011100;
#10000;
	data_in <= 24'b100110111000001001011101;
#10000;
	data_in <= 24'b100111001000001101011110;
#10000;
	data_in <= 24'b100111011000010001011111;
#10000;
	data_in <= 24'b100111011000010101100000;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b100111011000010001011110;
#10000;
	data_in <= 24'b100111101000010101011111;
#10000;
	data_in <= 24'b100111101000010101100000;
#10000;
	data_in <= 24'b100111111000011001100001;
#10000;
	data_in <= 24'b100111111000011001100010;
#10000;
	data_in <= 24'b101000001000100001100010;
#10000;
	data_in <= 24'b101000001000100101100011;
#10000;
	data_in <= 24'b101000001000011001100001;
#10000;
	data_in <= 24'b101000001000011101100010;
#10000;
	data_in <= 24'b101000011000100001100011;
#10000;
	data_in <= 24'b101000101000100101100100;
#10000;
	data_in <= 24'b101000111000101001100101;
#10000;
	data_in <= 24'b101000101000101001100110;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101001011000110101100111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010100111000001001011;
#10000;
	data_in <= 24'b100010100111000101001011;
#10000;
	data_in <= 24'b100010110111000101001011;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010100111001001001100;
#10000;
	data_in <= 24'b100011010111010001001110;
#10000;
	data_in <= 24'b100011010111010101001111;
#10000;
	data_in <= 24'b100011100111010101001111;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111011001010001;
#10000;
	data_in <= 24'b100100100111100101010011;
#10000;
	data_in <= 24'b100100100111100101010100;
#10000;
	data_in <= 24'b100100010111100001010100;
#10000;
	data_in <= 24'b100100010111100001010101;
#10000;
	data_in <= 24'b100100010111100101010101;
#10000;
	data_in <= 24'b100100010111100101010110;
#10000;
	data_in <= 24'b100100100111101001010101;
#10000;
	data_in <= 24'b100100100111101001010101;
#10000;
	data_in <= 24'b100101010111110001010111;
#10000;
	data_in <= 24'b100101010111110001010111;
#10000;
	data_in <= 24'b100101010111110001011000;
#10000;
	data_in <= 24'b100101100111110101011001;
#10000;
	data_in <= 24'b100101100111111001011001;
#10000;
	data_in <= 24'b100101100111111001011010;
#10000;
	data_in <= 24'b100101100111111001011010;
#10000;
	data_in <= 24'b100101110111111101011001;
#10000;
	data_in <= 24'b100110001000000001011100;
#10000;
	data_in <= 24'b100110011000000001011100;
#10000;
	data_in <= 24'b100110101000000101011100;
#10000;
	data_in <= 24'b100110111000000101011101;
#10000;
	data_in <= 24'b100110111000001101011101;
#10000;
	data_in <= 24'b100110111000001101011110;
#10000;
	data_in <= 24'b100110111000001101011110;
#10000;
	data_in <= 24'b100110101000001001011110;
#10000;
	data_in <= 24'b100111011000011001100001;
#10000;
	data_in <= 24'b100111101000011001100001;
#10000;
	data_in <= 24'b100111101000011001100001;
#10000;
	data_in <= 24'b100111011000011001100001;
#10000;
	data_in <= 24'b100111011000011001100001;
#10000;
	data_in <= 24'b100111011000011001100010;
#10000;
	data_in <= 24'b100111101000011001100010;
#10000;
	data_in <= 24'b100111111000011001100011;
#10000;
	data_in <= 24'b101000011000100101100100;
#10000;
	data_in <= 24'b101000011000100101100100;
#10000;
	data_in <= 24'b101000011000100101100100;
#10000;
	data_in <= 24'b101000011000101001100100;
#10000;
	data_in <= 24'b101000101000101001100101;
#10000;
	data_in <= 24'b101000101000101001100110;
#10000;
	data_in <= 24'b101000101000101001100110;
#10000;
	data_in <= 24'b101000101000101001100111;
#10000;
	data_in <= 24'b101001001000110001101000;
#10000;
	data_in <= 24'b101001011000110001101001;
#10000;
	data_in <= 24'b101001011000110001101001;
#10000;
	data_in <= 24'b101001001000110001101001;
#10000;
	data_in <= 24'b101001101000110101101010;
#10000;
	data_in <= 24'b101001111000111101101011;
#10000;
	data_in <= 24'b101001111000111101101011;
#10000;
	data_in <= 24'b101001011000110101101010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010110111001001001101;
#10000;
	data_in <= 24'b100011000111001001001110;
#10000;
	data_in <= 24'b100011000111001001001101;
#10000;
	data_in <= 24'b100011000111001101001101;
#10000;
	data_in <= 24'b100011000111001101001101;
#10000;
	data_in <= 24'b100010110111001101001110;
#10000;
	data_in <= 24'b100010110111001101001110;
#10000;
	data_in <= 24'b100010110111001101001110;
#10000;
	data_in <= 24'b100011100111011001010010;
#10000;
	data_in <= 24'b100011110111011001010010;
#10000;
	data_in <= 24'b100011110111011001010010;
#10000;
	data_in <= 24'b100011110111011101010010;
#10000;
	data_in <= 24'b100011110111011101010010;
#10000;
	data_in <= 24'b100011100111011101010011;
#10000;
	data_in <= 24'b100011100111011101010011;
#10000;
	data_in <= 24'b100011100111011101010011;
#10000;
	data_in <= 24'b100100110111101001010110;
#10000;
	data_in <= 24'b100101000111101001010111;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100100110111101101010110;
#10000;
	data_in <= 24'b100100110111101101010110;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100101110111111101011010;
#10000;
	data_in <= 24'b100110000111111101011010;
#10000;
	data_in <= 24'b100101110111111001011011;
#10000;
	data_in <= 24'b100110000111111101011011;
#10000;
	data_in <= 24'b100110001000000001011011;
#10000;
	data_in <= 24'b100101110111111101011100;
#10000;
	data_in <= 24'b100101110111111101011100;
#10000;
	data_in <= 24'b100101110111111101011100;
#10000;
	data_in <= 24'b100110111000001101011110;
#10000;
	data_in <= 24'b100110111000001101011111;
#10000;
	data_in <= 24'b100111001000001001011111;
#10000;
	data_in <= 24'b100110111000001101100000;
#10000;
	data_in <= 24'b100110111000010001100000;
#10000;
	data_in <= 24'b100110111000001101100001;
#10000;
	data_in <= 24'b100110111000010001100001;
#10000;
	data_in <= 24'b100111001000010001100001;
#10000;
	data_in <= 24'b100111101000011001100100;
#10000;
	data_in <= 24'b100111111000011001100011;
#10000;
	data_in <= 24'b101000001000011001100011;
#10000;
	data_in <= 24'b101000001000011101100011;
#10000;
	data_in <= 24'b101000001000100001100100;
#10000;
	data_in <= 24'b101000001000100001100111;
#10000;
	data_in <= 24'b101000001000100001100110;
#10000;
	data_in <= 24'b100111111000011101100011;
#10000;
	data_in <= 24'b101000101000101101100111;
#10000;
	data_in <= 24'b101000111000101101101000;
#10000;
	data_in <= 24'b101001001000101101101000;
#10000;
	data_in <= 24'b101000111000101101101000;
#10000;
	data_in <= 24'b101000011000100101100101;
#10000;
	data_in <= 24'b100111011000010001011111;
#10000;
	data_in <= 24'b100110101000001001011111;
#10000;
	data_in <= 24'b100110011000010101100110;
#10000;
	data_in <= 24'b101001011000111001101100;
#10000;
	data_in <= 24'b101001111000111101101101;
#10000;
	data_in <= 24'b101001001000101001100111;
#10000;
	data_in <= 24'b100111101000011001100011;
#10000;
	data_in <= 24'b100111001000101101101110;
#10000;
	data_in <= 24'b101000011001101110001011;
#10000;
	data_in <= 24'b101010001010110110101000;
#10000;
	data_in <= 24'b101011101011101010111100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010110111001101001110;
#10000;
	data_in <= 24'b100010110111001101001110;
#10000;
	data_in <= 24'b100010110111001101001110;
#10000;
	data_in <= 24'b100011000111001101001101;
#10000;
	data_in <= 24'b100011000111001101001101;
#10000;
	data_in <= 24'b100011000111001001001101;
#10000;
	data_in <= 24'b100011000111001001001110;
#10000;
	data_in <= 24'b100010110111001001001101;
#10000;
	data_in <= 24'b100011100111011101010011;
#10000;
	data_in <= 24'b100011100111011101010011;
#10000;
	data_in <= 24'b100011100111011101010011;
#10000;
	data_in <= 24'b100011110111011101010010;
#10000;
	data_in <= 24'b100011110111011101010010;
#10000;
	data_in <= 24'b100011110111011001010010;
#10000;
	data_in <= 24'b100011110111011001010010;
#10000;
	data_in <= 24'b100011100111011001010010;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100100110111101101010110;
#10000;
	data_in <= 24'b100100110111101101010110;
#10000;
	data_in <= 24'b100100110111101101010111;
#10000;
	data_in <= 24'b100101000111101001010111;
#10000;
	data_in <= 24'b100100110111101001010110;
#10000;
	data_in <= 24'b100101110111111101011100;
#10000;
	data_in <= 24'b100101110111111101011100;
#10000;
	data_in <= 24'b100101110111111101011100;
#10000;
	data_in <= 24'b100101111000000001011011;
#10000;
	data_in <= 24'b100101110111111101011011;
#10000;
	data_in <= 24'b100101110111111001011010;
#10000;
	data_in <= 24'b100110000111111001011010;
#10000;
	data_in <= 24'b100101110111111001011010;
#10000;
	data_in <= 24'b100111001000010101100010;
#10000;
	data_in <= 24'b100111001000010101100010;
#10000;
	data_in <= 24'b100111001000010101100011;
#10000;
	data_in <= 24'b100111001000010101100010;
#10000;
	data_in <= 24'b100111001000010101100010;
#10000;
	data_in <= 24'b100111001000010001100001;
#10000;
	data_in <= 24'b100111001000010001100001;
#10000;
	data_in <= 24'b100110111000001101011111;
#10000;
	data_in <= 24'b100111011000010001100000;
#10000;
	data_in <= 24'b100111001000001001011110;
#10000;
	data_in <= 24'b100110111000001001011101;
#10000;
	data_in <= 24'b100110111000000101011011;
#10000;
	data_in <= 24'b100110111000000101011011;
#10000;
	data_in <= 24'b100110111000000101011100;
#10000;
	data_in <= 24'b100111001000001001011110;
#10000;
	data_in <= 24'b100111011000010001100000;
#10000;
	data_in <= 24'b100110111000101001101111;
#10000;
	data_in <= 24'b100111001000111101111000;
#10000;
	data_in <= 24'b100111011001001001111101;
#10000;
	data_in <= 24'b100111011001010110000001;
#10000;
	data_in <= 24'b100111011001010001111111;
#10000;
	data_in <= 24'b100111011001000101111010;
#10000;
	data_in <= 24'b100110111000110101110100;
#10000;
	data_in <= 24'b100110011000011101101010;
#10000;
	data_in <= 24'b101100011100001011001000;
#10000;
	data_in <= 24'b101101001100011011001110;
#10000;
	data_in <= 24'b101101011100011111010001;
#10000;
	data_in <= 24'b101101011100100111010010;
#10000;
	data_in <= 24'b101101011100100011010010;
#10000;
	data_in <= 24'b101101011100011111010000;
#10000;
	data_in <= 24'b101100111100010011001011;
#10000;
	data_in <= 24'b101100001011111011000011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010100111001001001100;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010110111001001001100;
#10000;
	data_in <= 24'b100010110111000101001011;
#10000;
	data_in <= 24'b100010100111000101001011;
#10000;
	data_in <= 24'b100010100111000001001011;
#10000;
	data_in <= 24'b100011100111011001010001;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111011001010000;
#10000;
	data_in <= 24'b100011100111010101001111;
#10000;
	data_in <= 24'b100011010111010101001111;
#10000;
	data_in <= 24'b100011010111010001001110;
#10000;
	data_in <= 24'b100100100111101001010101;
#10000;
	data_in <= 24'b100100100111101001010101;
#10000;
	data_in <= 24'b100100010111100101010110;
#10000;
	data_in <= 24'b100100010111100101010101;
#10000;
	data_in <= 24'b100100010111100001010101;
#10000;
	data_in <= 24'b100100010111100001010100;
#10000;
	data_in <= 24'b100100100111100101010100;
#10000;
	data_in <= 24'b100100100111100101010011;
#10000;
	data_in <= 24'b100101100111111101011001;
#10000;
	data_in <= 24'b100101100111111001011010;
#10000;
	data_in <= 24'b100101100111111001011010;
#10000;
	data_in <= 24'b100101100111111001011001;
#10000;
	data_in <= 24'b100101100111110101011001;
#10000;
	data_in <= 24'b100101010111110001011000;
#10000;
	data_in <= 24'b100101010111110001010111;
#10000;
	data_in <= 24'b100101010111110001010111;
#10000;
	data_in <= 24'b100110111000001101011111;
#10000;
	data_in <= 24'b100110101000001001011110;
#10000;
	data_in <= 24'b100110101000001101011101;
#10000;
	data_in <= 24'b100110111000001101011101;
#10000;
	data_in <= 24'b100110111000000101011101;
#10000;
	data_in <= 24'b100110101000000101011100;
#10000;
	data_in <= 24'b100110011000000001011100;
#10000;
	data_in <= 24'b100110001000000001011100;
#10000;
	data_in <= 24'b100111111000011001100010;
#10000;
	data_in <= 24'b100111111000100001100100;
#10000;
	data_in <= 24'b100111101000011101100011;
#10000;
	data_in <= 24'b100111011000011101100010;
#10000;
	data_in <= 24'b100111011000011001100000;
#10000;
	data_in <= 24'b100111101000011001100001;
#10000;
	data_in <= 24'b100111101000011001100001;
#10000;
	data_in <= 24'b100111011000011001100001;
#10000;
	data_in <= 24'b100110011000001001100000;
#10000;
	data_in <= 24'b100110101000000101011100;
#10000;
	data_in <= 24'b100111111000010101100000;
#10000;
	data_in <= 24'b101000101000101001100101;
#10000;
	data_in <= 24'b101000101000101001100110;
#10000;
	data_in <= 24'b101000011000101001100101;
#10000;
	data_in <= 24'b101000011000100101100100;
#10000;
	data_in <= 24'b101000011000100101100100;
#10000;
	data_in <= 24'b101010111011010110110100;
#10000;
	data_in <= 24'b101001011010010110011011;
#10000;
	data_in <= 24'b100111011001001001111100;
#10000;
	data_in <= 24'b100110111000011001100101;
#10000;
	data_in <= 24'b101000001000011001100010;
#10000;
	data_in <= 24'b101001001000110001101000;
#10000;
	data_in <= 24'b101001011000110101101010;
#10000;
	data_in <= 24'b101000111000110001101000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010100111000101001011;
#10000;
	data_in <= 24'b100010100111000001001011;
#10000;
	data_in <= 24'b100010100111000001001001;
#10000;
	data_in <= 24'b100010010110111101001001;
#10000;
	data_in <= 24'b100010000110111001000111;
#10000;
	data_in <= 24'b100010000110111001000110;
#10000;
	data_in <= 24'b100001110110110101000110;
#10000;
	data_in <= 24'b100001100110110001000101;
#10000;
	data_in <= 24'b100011010111010101001110;
#10000;
	data_in <= 24'b100011010111010001001110;
#10000;
	data_in <= 24'b100011000111010001001101;
#10000;
	data_in <= 24'b100010110111001101001101;
#10000;
	data_in <= 24'b100010110111001001001011;
#10000;
	data_in <= 24'b100010110111000101001010;
#10000;
	data_in <= 24'b100010110111000101001010;
#10000;
	data_in <= 24'b100010100111000001001001;
#10000;
	data_in <= 24'b100100010111100001010011;
#10000;
	data_in <= 24'b100100010111100001010010;
#10000;
	data_in <= 24'b100100000111011101010010;
#10000;
	data_in <= 24'b100100000111011101010001;
#10000;
	data_in <= 24'b100011110111011001001111;
#10000;
	data_in <= 24'b100011100111010101001111;
#10000;
	data_in <= 24'b100011100111010001001110;
#10000;
	data_in <= 24'b100011010111001101001101;
#10000;
	data_in <= 24'b100101010111110001010111;
#10000;
	data_in <= 24'b100101000111101101010101;
#10000;
	data_in <= 24'b100101000111101101010101;
#10000;
	data_in <= 24'b100100110111101001010100;
#10000;
	data_in <= 24'b100100110111101001010100;
#10000;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b100100010111100001010001;
#10000;
	data_in <= 24'b100110011000000001011100;
#10000;
	data_in <= 24'b100110011000000001011011;
#10000;
	data_in <= 24'b100101110111111001011010;
#10000;
	data_in <= 24'b100101100111110101011001;
#10000;
	data_in <= 24'b100101100111110101011000;
#10000;
	data_in <= 24'b100101100111110101010111;
#10000;
	data_in <= 24'b100101010111110001010110;
#10000;
	data_in <= 24'b100101010111101101010101;
#10000;
	data_in <= 24'b100111011000010101100000;
#10000;
	data_in <= 24'b100111011000010001011111;
#10000;
	data_in <= 24'b100111001000001101011110;
#10000;
	data_in <= 24'b100110111000001001011101;
#10000;
	data_in <= 24'b100110111000001001011100;
#10000;
	data_in <= 24'b100110101000000101011100;
#10000;
	data_in <= 24'b100110101000000101011011;
#10000;
	data_in <= 24'b100110011000000001011010;
#10000;
	data_in <= 24'b101000001000100001100011;
#10000;
	data_in <= 24'b100111111000011101100010;
#10000;
	data_in <= 24'b100111111000011001100010;
#10000;
	data_in <= 24'b100111101000010101100001;
#10000;
	data_in <= 24'b100111101000010101100000;
#10000;
	data_in <= 24'b100111101000010101011111;
#10000;
	data_in <= 24'b100111011000010001011110;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101001011000110001100111;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101000101000101001100101;
#10000;
	data_in <= 24'b101000001000100001100100;
#10000;
	data_in <= 24'b101000011000100001100011;
#10000;
	data_in <= 24'b101000001000011101100010;
#10000;
	data_in <= 24'b101000001000011001100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100001100110110001000011;
#10000;
	data_in <= 24'b100001010110101001000010;
#10000;
	data_in <= 24'b100001010110100001000010;
#10000;
	data_in <= 24'b100001000110100001000000;
#10000;
	data_in <= 24'b100000100110011100111111;
#10000;
	data_in <= 24'b100000010110011100111110;
#10000;
	data_in <= 24'b011111110110010100111101;
#10000;
	data_in <= 24'b011111110110010000111011;
#10000;
	data_in <= 24'b100010010110111101001000;
#10000;
	data_in <= 24'b100010010110111001000110;
#10000;
	data_in <= 24'b100010000110110101000101;
#10000;
	data_in <= 24'b100010000110110001000101;
#10000;
	data_in <= 24'b100001110110101101000100;
#10000;
	data_in <= 24'b100001000110101001000010;
#10000;
	data_in <= 24'b100000110110100101000000;
#10000;
	data_in <= 24'b100000100110011100111111;
#10000;
	data_in <= 24'b100011010111001001001100;
#10000;
	data_in <= 24'b100011000111000101001010;
#10000;
	data_in <= 24'b100010110111000001001001;
#10000;
	data_in <= 24'b100010110110111101001001;
#10000;
	data_in <= 24'b100010100110111001001000;
#10000;
	data_in <= 24'b100010000110110101000110;
#10000;
	data_in <= 24'b100001100110101101000100;
#10000;
	data_in <= 24'b100001010110101001000010;
#10000;
	data_in <= 24'b100100000111011001010000;
#10000;
	data_in <= 24'b100100000111010101001110;
#10000;
	data_in <= 24'b100011110111010001001101;
#10000;
	data_in <= 24'b100011100111001101001100;
#10000;
	data_in <= 24'b100011000111001001001010;
#10000;
	data_in <= 24'b100011000111000001001001;
#10000;
	data_in <= 24'b100010100110111001001000;
#10000;
	data_in <= 24'b100010010110111001000110;
#10000;
	data_in <= 24'b100101000111101001010100;
#10000;
	data_in <= 24'b100100110111100001010011;
#10000;
	data_in <= 24'b100100110111100001010010;
#10000;
	data_in <= 24'b100100100111011101010000;
#10000;
	data_in <= 24'b100100000111011001001110;
#10000;
	data_in <= 24'b100011110111010101001110;
#10000;
	data_in <= 24'b100011100111001001001100;
#10000;
	data_in <= 24'b100011010111000101001010;
#10000;
	data_in <= 24'b100110000111110101010111;
#10000;
	data_in <= 24'b100101110111110001010110;
#10000;
	data_in <= 24'b100101110111110001010110;
#10000;
	data_in <= 24'b100101100111101101010100;
#10000;
	data_in <= 24'b100101000111101001010010;
#10000;
	data_in <= 24'b100100100111100101010001;
#10000;
	data_in <= 24'b100100010111011101010000;
#10000;
	data_in <= 24'b100100000111010101001110;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100110111000000001011010;
#10000;
	data_in <= 24'b100110100111111101011001;
#10000;
	data_in <= 24'b100110010111111001010111;
#10000;
	data_in <= 24'b100110000111110101010110;
#10000;
	data_in <= 24'b100101100111101101010100;
#10000;
	data_in <= 24'b100101000111101001010011;
#10000;
	data_in <= 24'b100100100111100101010001;
#10000;
	data_in <= 24'b100111111000010101011111;
#10000;
	data_in <= 24'b100111101000010001011110;
#10000;
	data_in <= 24'b100111101000001101011101;
#10000;
	data_in <= 24'b100111001000001001011100;
#10000;
	data_in <= 24'b100110101000000001011010;
#10000;
	data_in <= 24'b100110100111111101011001;
#10000;
	data_in <= 24'b100110000111110101010111;
#10000;
	data_in <= 24'b100101100111110001010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011111100110001100111001;
#10000;
	data_in <= 24'b011111010110000100111000;
#10000;
	data_in <= 24'b011111000110000000110111;
#10000;
	data_in <= 24'b011110110101111100110101;
#10000;
	data_in <= 24'b011110100101111000110011;
#10000;
	data_in <= 24'b011110000101110000110001;
#10000;
	data_in <= 24'b011101110101100100101111;
#10000;
	data_in <= 24'b011101100101100000101111;
#10000;
	data_in <= 24'b100000010110011000111101;
#10000;
	data_in <= 24'b100000000110010100111011;
#10000;
	data_in <= 24'b011111110110001100111011;
#10000;
	data_in <= 24'b011111100110001000111001;
#10000;
	data_in <= 24'b011111010110000000110110;
#10000;
	data_in <= 24'b011111000101111000110101;
#10000;
	data_in <= 24'b011110100101110100110011;
#10000;
	data_in <= 24'b011110000101101100110010;
#10000;
	data_in <= 24'b100001010110100101000001;
#10000;
	data_in <= 24'b100000110110100000111111;
#10000;
	data_in <= 24'b100000100110011000111110;
#10000;
	data_in <= 24'b100000000110010000111100;
#10000;
	data_in <= 24'b100000000110001100111010;
#10000;
	data_in <= 24'b011111100110001000111001;
#10000;
	data_in <= 24'b011111000110000000110111;
#10000;
	data_in <= 24'b011110100101111000110100;
#10000;
	data_in <= 24'b100001110110110001000100;
#10000;
	data_in <= 24'b100001100110101101000011;
#10000;
	data_in <= 24'b100001010110101001000001;
#10000;
	data_in <= 24'b100001000110100000111111;
#10000;
	data_in <= 24'b100000110110010100111101;
#10000;
	data_in <= 24'b100000010110010100111011;
#10000;
	data_in <= 24'b011111110110001100111010;
#10000;
	data_in <= 24'b011111100110000100110111;
#10000;
	data_in <= 24'b100010110111000001001000;
#10000;
	data_in <= 24'b100010100110111101000111;
#10000;
	data_in <= 24'b100010000110110101000101;
#10000;
	data_in <= 24'b100001110110101101000011;
#10000;
	data_in <= 24'b100001100110100101000001;
#10000;
	data_in <= 24'b100001000110011100111111;
#10000;
	data_in <= 24'b100000100110011000111101;
#10000;
	data_in <= 24'b100000000110010000111010;
#10000;
	data_in <= 24'b100011100111001101001100;
#10000;
	data_in <= 24'b100011010111001001001010;
#10000;
	data_in <= 24'b100011000111000101001000;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100010010110110001000100;
#10000;
	data_in <= 24'b100010000110101101000011;
#10000;
	data_in <= 24'b100001100110100101000000;
#10000;
	data_in <= 24'b100000110110011100111101;
#10000;
	data_in <= 24'b100100100111011101001111;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b100011110111010001001011;
#10000;
	data_in <= 24'b100011010111001001001000;
#10000;
	data_in <= 24'b100011000110111101000111;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100010000110110001000010;
#10000;
	data_in <= 24'b100001100110101001000000;
#10000;
	data_in <= 24'b100101010111101001010011;
#10000;
	data_in <= 24'b100101000111100001010000;
#10000;
	data_in <= 24'b100100100111011101001111;
#10000;
	data_in <= 24'b100100000111010101001101;
#10000;
	data_in <= 24'b100011100111001001001010;
#10000;
	data_in <= 24'b100011000111000001001001;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100010000110110001000011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011101000101011100101100;
#10000;
	data_in <= 24'b011100100101011000101010;
#10000;
	data_in <= 24'b011100010101010000101001;
#10000;
	data_in <= 24'b011011110101000100100111;
#10000;
	data_in <= 24'b011011010100111100100100;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011010100100110000100000;
#10000;
	data_in <= 24'b011010010100101000011110;
#10000;
	data_in <= 24'b011101100101100100110000;
#10000;
	data_in <= 24'b011101000101100000101101;
#10000;
	data_in <= 24'b011100110101011100101011;
#10000;
	data_in <= 24'b011100010101010000101010;
#10000;
	data_in <= 24'b011100000101001000100111;
#10000;
	data_in <= 24'b011011100101000000100101;
#10000;
	data_in <= 24'b011011000100111000100011;
#10000;
	data_in <= 24'b011010110100110000100000;
#10000;
	data_in <= 24'b011110010101110000110010;
#10000;
	data_in <= 24'b011101110101101000110000;
#10000;
	data_in <= 24'b011101010101100100101110;
#10000;
	data_in <= 24'b011101000101011100101100;
#10000;
	data_in <= 24'b011100100101010000101001;
#10000;
	data_in <= 24'b011100000101001000100111;
#10000;
	data_in <= 24'b011011110101000000100101;
#10000;
	data_in <= 24'b011011010100111000100011;
#10000;
	data_in <= 24'b011111000101111100110101;
#10000;
	data_in <= 24'b011110100101110100110011;
#10000;
	data_in <= 24'b011110000101101100110001;
#10000;
	data_in <= 24'b011101100101100100101110;
#10000;
	data_in <= 24'b011101000101011000101011;
#10000;
	data_in <= 24'b011100100101010000101001;
#10000;
	data_in <= 24'b011100000101001100100111;
#10000;
	data_in <= 24'b011011110101000000100101;
#10000;
	data_in <= 24'b011111100110001000111000;
#10000;
	data_in <= 24'b011111010110000000110111;
#10000;
	data_in <= 24'b011110110101110100110011;
#10000;
	data_in <= 24'b011110000101101100110000;
#10000;
	data_in <= 24'b011101100101100100101111;
#10000;
	data_in <= 24'b011101010101011100101100;
#10000;
	data_in <= 24'b011100110101010100101010;
#10000;
	data_in <= 24'b011100010101001100101000;
#10000;
	data_in <= 24'b100000100110010100111011;
#10000;
	data_in <= 24'b100000000110001000111001;
#10000;
	data_in <= 24'b011111010110000000110110;
#10000;
	data_in <= 24'b011111000101111000110100;
#10000;
	data_in <= 24'b011110100101110000110010;
#10000;
	data_in <= 24'b011101110101100100101111;
#10000;
	data_in <= 24'b011101010101011100101100;
#10000;
	data_in <= 24'b011100110101010100101010;
#10000;
	data_in <= 24'b100001010110100000111110;
#10000;
	data_in <= 24'b100000100110010100111010;
#10000;
	data_in <= 24'b100000000110001000111001;
#10000;
	data_in <= 24'b011111010110000100110110;
#10000;
	data_in <= 24'b011111000101111100110100;
#10000;
	data_in <= 24'b011110100101110000110000;
#10000;
	data_in <= 24'b011101110101100100101101;
#10000;
	data_in <= 24'b011101010101011100101011;
#10000;
	data_in <= 24'b100001110110101001000010;
#10000;
	data_in <= 24'b100001010110011100111110;
#10000;
	data_in <= 24'b100000100110010000111011;
#10000;
	data_in <= 24'b100000000110001100111010;
#10000;
	data_in <= 24'b011111100110000000110111;
#10000;
	data_in <= 24'b011111000101111000110100;
#10000;
	data_in <= 24'b011110010101101100110001;
#10000;
	data_in <= 24'b011101110101100100101110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011110000101101000110001;
#10000;
	data_in <= 24'b011110110101110100110011;
#10000;
	data_in <= 24'b011111010101111100110110;
#10000;
	data_in <= 24'b011111110110001000111001;
#10000;
	data_in <= 24'b100000100110010100111100;
#10000;
	data_in <= 24'b100001010110011100111110;
#10000;
	data_in <= 24'b100001110110101001000001;
#10000;
	data_in <= 24'b100010010110110001000100;
#10000;
	data_in <= 24'b011110100101110100110010;
#10000;
	data_in <= 24'b011111010101111100110101;
#10000;
	data_in <= 24'b011111110110001000111000;
#10000;
	data_in <= 24'b100000010110010100111011;
#10000;
	data_in <= 24'b100001000110011100111110;
#10000;
	data_in <= 24'b100001110110101001000001;
#10000;
	data_in <= 24'b100010010110110001000011;
#10000;
	data_in <= 24'b100010110110111101000110;
#10000;
	data_in <= 24'b011111000110000000110100;
#10000;
	data_in <= 24'b011111100110000100110111;
#10000;
	data_in <= 24'b100000000110010000111010;
#10000;
	data_in <= 24'b100000110110011100111110;
#10000;
	data_in <= 24'b100001110110101001000001;
#10000;
	data_in <= 24'b100010010110110001000011;
#10000;
	data_in <= 24'b100010110110111001000101;
#10000;
	data_in <= 24'b100011100111001001001001;
#10000;
	data_in <= 24'b011111010110000000110101;
#10000;
	data_in <= 24'b100000000110001100111001;
#10000;
	data_in <= 24'b100000110110011100111100;
#10000;
	data_in <= 24'b100001100110100101000000;
#10000;
	data_in <= 24'b100010000110101101000010;
#10000;
	data_in <= 24'b100010110110111001000101;
#10000;
	data_in <= 24'b100011010111000101001000;
#10000;
	data_in <= 24'b100011110111010001001011;
#10000;
	data_in <= 24'b011111100110000100111000;
#10000;
	data_in <= 24'b100000010110010000111011;
#10000;
	data_in <= 24'b100001000110100000111111;
#10000;
	data_in <= 24'b100001110110101101000010;
#10000;
	data_in <= 24'b100010100110110101000101;
#10000;
	data_in <= 24'b100011010111000001000111;
#10000;
	data_in <= 24'b100011110111001101001011;
#10000;
	data_in <= 24'b100100010111010101001101;
#10000;
	data_in <= 24'b011111110110001100111001;
#10000;
	data_in <= 24'b100000100110011000111101;
#10000;
	data_in <= 24'b100001010110101001000000;
#10000;
	data_in <= 24'b100010000110110101000011;
#10000;
	data_in <= 24'b100011000111000001000111;
#10000;
	data_in <= 24'b100011110111001101001010;
#10000;
	data_in <= 24'b100100010111011001001101;
#10000;
	data_in <= 24'b100100110111100001001111;
#10000;
	data_in <= 24'b100000010110010000111011;
#10000;
	data_in <= 24'b100001000110100000111110;
#10000;
	data_in <= 24'b100001110110110001000001;
#10000;
	data_in <= 24'b100010110110111001000101;
#10000;
	data_in <= 24'b100011110111001001001001;
#10000;
	data_in <= 24'b100100000111010101001100;
#10000;
	data_in <= 24'b100100110111011101001111;
#10000;
	data_in <= 24'b100101010111101001010010;
#10000;
	data_in <= 24'b100001000110011000111101;
#10000;
	data_in <= 24'b100001110110101001000000;
#10000;
	data_in <= 24'b100010010110110101000011;
#10000;
	data_in <= 24'b100011010111000001000111;
#10000;
	data_in <= 24'b100100010111010001001011;
#10000;
	data_in <= 24'b100100110111011001001110;
#10000;
	data_in <= 24'b100101010111100101010001;
#10000;
	data_in <= 24'b100110000111110001010100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100011000111000001001000;
#10000;
	data_in <= 24'b100011100111001101001100;
#10000;
	data_in <= 24'b100100010111010101001101;
#10000;
	data_in <= 24'b100100100111011101001111;
#10000;
	data_in <= 24'b100101000111100101010001;
#10000;
	data_in <= 24'b100101100111101101010011;
#10000;
	data_in <= 24'b100101110111110101010110;
#10000;
	data_in <= 24'b100011010111001001001000;
#10000;
	data_in <= 24'b100011110111010001001011;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b100100110111100001010000;
#10000;
	data_in <= 24'b100101010111101001010011;
#10000;
	data_in <= 24'b100101110111110101010100;
#10000;
	data_in <= 24'b100110010111111001010111;
#10000;
	data_in <= 24'b100110101000000001011010;
#10000;
	data_in <= 24'b100100000111010001001100;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b100100110111100101010001;
#10000;
	data_in <= 24'b100101010111101101010100;
#10000;
	data_in <= 24'b100110000111110101010110;
#10000;
	data_in <= 24'b100110100111111101011000;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b100100110111100101010000;
#10000;
	data_in <= 24'b100101010111101101010011;
#10000;
	data_in <= 24'b100101110111110101010110;
#10000;
	data_in <= 24'b100110100111111101011000;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100111101000010001011101;
#10000;
	data_in <= 24'b101000001000011001011111;
#10000;
	data_in <= 24'b100100110111100001010001;
#10000;
	data_in <= 24'b100101010111101101010011;
#10000;
	data_in <= 24'b100110000111111001010110;
#10000;
	data_in <= 24'b100110101000000001011001;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100111101000001101011101;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b101000111000100101100010;
#10000;
	data_in <= 24'b100101010111101001010011;
#10000;
	data_in <= 24'b100110000111111001010110;
#10000;
	data_in <= 24'b100110101000000001011001;
#10000;
	data_in <= 24'b100111001000001001011011;
#10000;
	data_in <= 24'b100111011000010001011101;
#10000;
	data_in <= 24'b101000011000011101100000;
#10000;
	data_in <= 24'b101000111000101001100011;
#10000;
	data_in <= 24'b101001011000110001100101;
#10000;
	data_in <= 24'b100110000111110101010110;
#10000;
	data_in <= 24'b100110101000000001011000;
#10000;
	data_in <= 24'b100111001000001101011011;
#10000;
	data_in <= 24'b100111101000010101011101;
#10000;
	data_in <= 24'b101000001000011101100000;
#10000;
	data_in <= 24'b101000111000101001100010;
#10000;
	data_in <= 24'b101001101000110101100101;
#10000;
	data_in <= 24'b101001111000111001100111;
#10000;
	data_in <= 24'b100110100111111001011000;
#10000;
	data_in <= 24'b100111011000000101011011;
#10000;
	data_in <= 24'b100111101000010001011101;
#10000;
	data_in <= 24'b101000011000011101100001;
#10000;
	data_in <= 24'b101001001000100101100011;
#10000;
	data_in <= 24'b101001111000110001100110;
#10000;
	data_in <= 24'b101010001000111001100111;
#10000;
	data_in <= 24'b101010101001000001101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100110010111111101011000;
#10000;
	data_in <= 24'b100110111000000001011010;
#10000;
	data_in <= 24'b100111011000000101011101;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b100111111000010001011111;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b101000011000011101100001;
#10000;
	data_in <= 24'b101000101000100001100011;
#10000;
	data_in <= 24'b100111001000001001011011;
#10000;
	data_in <= 24'b100111101000001101011101;
#10000;
	data_in <= 24'b100111111000010101011111;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b101000101000100101100010;
#10000;
	data_in <= 24'b101001001000101101100100;
#10000;
	data_in <= 24'b101001011000101101100110;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
	data_in <= 24'b100111111000010101011110;
#10000;
	data_in <= 24'b101000001000011101100000;
#10000;
	data_in <= 24'b101000101000100001100011;
#10000;
	data_in <= 24'b101000111000101001100100;
#10000;
	data_in <= 24'b101001011000110101100110;
#10000;
	data_in <= 24'b101001101000111001101000;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101000101000100001100001;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b101001001000101101100101;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101001111000111101101000;
#10000;
	data_in <= 24'b101010001001000001101010;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101010111001001001101101;
#10000;
	data_in <= 24'b101001001000101001100100;
#10000;
	data_in <= 24'b101001101000110001100111;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101010001001000101101010;
#10000;
	data_in <= 24'b101010011001001001101100;
#10000;
	data_in <= 24'b101010111001001101101110;
#10000;
	data_in <= 24'b101011011001010001110000;
#10000;
	data_in <= 24'b101011101001010101110000;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101010001000111001101010;
#10000;
	data_in <= 24'b101010011001000001101011;
#10000;
	data_in <= 24'b101010111001010001101110;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b101011101001011001110001;
#10000;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b101010011001000001101001;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101011001001010001101110;
#10000;
	data_in <= 24'b101011101001011001110000;
#10000;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b101100101001101001110101;
#10000;
	data_in <= 24'b101100111001101101110110;
#10000;
	data_in <= 24'b101011001001001001101101;
#10000;
	data_in <= 24'b101011101001010001101111;
#10000;
	data_in <= 24'b101011111001011001110001;
#10000;
	data_in <= 24'b101100011001100001110010;
#10000;
	data_in <= 24'b101100101001101001110101;
#10000;
	data_in <= 24'b101100111001101101110110;
#10000;
	data_in <= 24'b101101011001110001111000;
#10000;
	data_in <= 24'b101101111001111001111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000111000100101100100;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101001011000110101101000;
#10000;
	data_in <= 24'b101001011000110101101001;
#10000;
	data_in <= 24'b101001101000111001101010;
#10000;
	data_in <= 24'b101001111000111101101010;
#10000;
	data_in <= 24'b101001111001000001101010;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101001111000111101101010;
#10000;
	data_in <= 24'b101010001001000001101011;
#10000;
	data_in <= 24'b101010011001000101101100;
#10000;
	data_in <= 24'b101010011001000101101101;
#10000;
	data_in <= 24'b101010101001001001101110;
#10000;
	data_in <= 24'b101011001001010001101111;
#10000;
	data_in <= 24'b101010011001000001101011;
#10000;
	data_in <= 24'b101010101001000101101101;
#10000;
	data_in <= 24'b101010111001001101101110;
#10000;
	data_in <= 24'b101011001001010001101111;
#10000;
	data_in <= 24'b101011001001010101110000;
#10000;
	data_in <= 24'b101011001001010101110010;
#10000;
	data_in <= 24'b101011101001011001110011;
#10000;
	data_in <= 24'b101011011001011001110010;
#10000;
	data_in <= 24'b101011001001001101101111;
#10000;
	data_in <= 24'b101011011001010001110000;
#10000;
	data_in <= 24'b101011011001011001110001;
#10000;
	data_in <= 24'b101011101001011101110010;
#10000;
	data_in <= 24'b101011111001100001110011;
#10000;
	data_in <= 24'b101100011001100101110101;
#10000;
	data_in <= 24'b101011111001100001110101;
#10000;
	data_in <= 24'b101100111001101101110110;
#10000;
	data_in <= 24'b101011111001010101110010;
#10000;
	data_in <= 24'b101100001001011101110100;
#10000;
	data_in <= 24'b101100001001100101110101;
#10000;
	data_in <= 24'b101100011001101001110101;
#10000;
	data_in <= 24'b101100111001101001110110;
#10000;
	data_in <= 24'b101100101001101001111000;
#10000;
	data_in <= 24'b101101001001110001111001;
#10000;
	data_in <= 24'b101001001001000001110001;
#10000;
	data_in <= 24'b101100011001100101110100;
#10000;
	data_in <= 24'b101100101001110001110111;
#10000;
	data_in <= 24'b101100111001110101111000;
#10000;
	data_in <= 24'b101101011001110101111000;
#10000;
	data_in <= 24'b101101011001111001111001;
#10000;
	data_in <= 24'b101101001001111001111011;
#10000;
	data_in <= 24'b101101111010000001111100;
#10000;
	data_in <= 24'b010111010101110101010101;
#10000;
	data_in <= 24'b101101001001110101111000;
#10000;
	data_in <= 24'b101101101001111101111010;
#10000;
	data_in <= 24'b101101111010000001111011;
#10000;
	data_in <= 24'b101110001010000001111100;
#10000;
	data_in <= 24'b101101111010000001111100;
#10000;
	data_in <= 24'b101111001010010010000000;
#10000;
	data_in <= 24'b100101111000100001101110;
#10000;
	data_in <= 24'b000110010010110000110111;
#10000;
	data_in <= 24'b101101111001111101111011;
#10000;
	data_in <= 24'b101110011010000101111101;
#10000;
	data_in <= 24'b101110101010001001111110;
#10000;
	data_in <= 24'b101110111010001101111111;
#10000;
	data_in <= 24'b101110101010001010000000;
#10000;
	data_in <= 24'b101111111010011010000010;
#10000;
	data_in <= 24'b010111010101110001010011;
#10000;
	data_in <= 24'b000000000001011000100111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101010001001000001101100;
#10000;
	data_in <= 24'b101010001000111101101100;
#10000;
	data_in <= 24'b101010011001000001101101;
#10000;
	data_in <= 24'b101010111001000001101100;
#10000;
	data_in <= 24'b101000101000101101101001;
#10000;
	data_in <= 24'b100110101000011101101001;
#10000;
	data_in <= 24'b100111011000100001101001;
#10000;
	data_in <= 24'b101010011001000101101110;
#10000;
	data_in <= 24'b101010111001001101101111;
#10000;
	data_in <= 24'b101011011001010001110000;
#10000;
	data_in <= 24'b101000101000110001101100;
#10000;
	data_in <= 24'b011110110111010101100101;
#10000;
	data_in <= 24'b010111100110010101100100;
#10000;
	data_in <= 24'b010100100101111001100011;
#10000;
	data_in <= 24'b010100100101110101100001;
#10000;
	data_in <= 24'b011001000110010001011011;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b100101101000011001101011;
#10000;
	data_in <= 24'b010100110101101101011100;
#10000;
	data_in <= 24'b001110110100111101011101;
#10000;
	data_in <= 24'b001111010101001101100001;
#10000;
	data_in <= 24'b010000000101011001100011;
#10000;
	data_in <= 24'b001100010100011101010101;
#10000;
	data_in <= 24'b001100000100010101010011;
#10000;
	data_in <= 24'b100101011000010101101011;
#10000;
	data_in <= 24'b001111100100101101010010;
#10000;
	data_in <= 24'b001011100100010001010100;
#10000;
	data_in <= 24'b001110100100111001011011;
#10000;
	data_in <= 24'b001111010101001001011111;
#10000;
	data_in <= 24'b001100100100100001010101;
#10000;
	data_in <= 24'b001101010100101001010111;
#10000;
	data_in <= 24'b100011011010000010101010;
#10000;
	data_in <= 24'b001111100100100101001101;
#10000;
	data_in <= 24'b001000010011100001001000;
#10000;
	data_in <= 24'b001011110100010101010001;
#10000;
	data_in <= 24'b001100000100011001010100;
#10000;
	data_in <= 24'b001010010100000101001111;
#10000;
	data_in <= 24'b001001010011110001001001;
#10000;
	data_in <= 24'b100000101001011110100010;
#10000;
	data_in <= 24'b101100101100011011010000;
#10000;
	data_in <= 24'b000100100010101000111010;
#10000;
	data_in <= 24'b001000110011100101000110;
#10000;
	data_in <= 24'b001000110011101001001000;
#10000;
	data_in <= 24'b001000010011100101000111;
#10000;
	data_in <= 24'b000100110010101000111001;
#10000;
	data_in <= 24'b011000110111100110000101;
#10000;
	data_in <= 24'b101100001100010011001110;
#10000;
	data_in <= 24'b101001101011101111000101;
#10000;
	data_in <= 24'b000100100010100100111000;
#10000;
	data_in <= 24'b000110010011000000111111;
#10000;
	data_in <= 24'b000110010011000101000000;
#10000;
	data_in <= 24'b000010100010001100110001;
#10000;
	data_in <= 24'b001100000100100001010101;
#10000;
	data_in <= 24'b101000111011100011000010;
#10000;
	data_in <= 24'b101001111011110011000110;
#10000;
	data_in <= 24'b101001111011110011000110;
#10000;
	data_in <= 24'b000011110010011100110101;
#10000;
	data_in <= 24'b000011110010011100110111;
#10000;
	data_in <= 24'b000010110010011000110101;
#10000;
	data_in <= 24'b000001010001110100101101;
#10000;
	data_in <= 24'b011110001000111010011001;
#10000;
	data_in <= 24'b101010101011111111001010;
#10000;
	data_in <= 24'b101001011011101011000100;
#10000;
	data_in <= 24'b101010001011111011001000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101010011001000101101110;
#10000;
	data_in <= 24'b101000011000100101100110;
#10000;
	data_in <= 24'b100111111000111101110110;
#10000;
	data_in <= 24'b101001011010011110011111;
#10000;
	data_in <= 24'b101011111011111111000101;
#10000;
	data_in <= 24'b101101001100100111010011;
#10000;
	data_in <= 24'b101101101100101011010110;
#10000;
	data_in <= 24'b101101101100101011010101;
#10000;
	data_in <= 24'b100011100111111101100101;
#10000;
	data_in <= 24'b101000111010001010010110;
#10000;
	data_in <= 24'b101011001011111011000101;
#10000;
	data_in <= 24'b101100111100100111010101;
#10000;
	data_in <= 24'b101100111100011111010001;
#10000;
	data_in <= 24'b101100101100010111001110;
#10000;
	data_in <= 24'b101100101100010111001110;
#10000;
	data_in <= 24'b101100011100010111001110;
#10000;
	data_in <= 24'b100011001001110110100011;
#10000;
	data_in <= 24'b101100111100011111010010;
#10000;
	data_in <= 24'b101011111100010011001111;
#10000;
	data_in <= 24'b101100001100001111001100;
#10000;
	data_in <= 24'b101011111100001111001101;
#10000;
	data_in <= 24'b101011111100001111001100;
#10000;
	data_in <= 24'b101011101100001111001100;
#10000;
	data_in <= 24'b101011011100001011001100;
#10000;
	data_in <= 24'b101100011100011011010001;
#10000;
	data_in <= 24'b101011001100000011001001;
#10000;
	data_in <= 24'b101011011100000111001010;
#10000;
	data_in <= 24'b101011011100001011001100;
#10000;
	data_in <= 24'b101011011100000111001011;
#10000;
	data_in <= 24'b101010111100000011001010;
#10000;
	data_in <= 24'b101010101011111111001010;
#10000;
	data_in <= 24'b101010011011111011001001;
#10000;
	data_in <= 24'b101010101011110111000111;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101010111100000111001010;
#10000;
	data_in <= 24'b101010111100000011001010;
#10000;
	data_in <= 24'b101010011011111011001000;
#10000;
	data_in <= 24'b101010001011110111001000;
#10000;
	data_in <= 24'b101001101011110011000111;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101010111100000011001010;
#10000;
	data_in <= 24'b101010101100000011001010;
#10000;
	data_in <= 24'b101010001011111011001000;
#10000;
	data_in <= 24'b101001111011110011000111;
#10000;
	data_in <= 24'b101001111011110011000111;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
	data_in <= 24'b101010101011111111001001;
#10000;
	data_in <= 24'b101001101011110111000111;
#10000;
	data_in <= 24'b101000101011101011000101;
#10000;
	data_in <= 24'b101000101011101011000100;
#10000;
	data_in <= 24'b101000011011100011000011;
#10000;
	data_in <= 24'b100111101011011111000010;
#10000;
	data_in <= 24'b101000011011100111000100;
#10000;
	data_in <= 24'b101001001011101111000101;
#10000;
	data_in <= 24'b101001001011110011000110;
#10000;
	data_in <= 24'b101100011100001111001011;
#10000;
	data_in <= 24'b110001111101001011010111;
#10000;
	data_in <= 24'b110100111101101111011111;
#10000;
	data_in <= 24'b110100101101101011011111;
#10000;
	data_in <= 24'b110000101100111111010101;
#10000;
	data_in <= 24'b101010001011110111000110;
#10000;
	data_in <= 24'b100111111011011111000011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101101101100101011010100;
#10000;
	data_in <= 24'b101101011100100111010011;
#10000;
	data_in <= 24'b101101011100100011010001;
#10000;
	data_in <= 24'b101101011100100011010001;
#10000;
	data_in <= 24'b101101011100100011010001;
#10000;
	data_in <= 24'b101101011100100011010010;
#10000;
	data_in <= 24'b101101101100100111010011;
#10000;
	data_in <= 24'b101101101100101011010100;
#10000;
	data_in <= 24'b101100011100010011001110;
#10000;
	data_in <= 24'b101100001100010011001101;
#10000;
	data_in <= 24'b101100001100010011001101;
#10000;
	data_in <= 24'b101100001100010011001110;
#10000;
	data_in <= 24'b101100001100010011001110;
#10000;
	data_in <= 24'b101100001100010011001101;
#10000;
	data_in <= 24'b101100011100010111001101;
#10000;
	data_in <= 24'b101100011100010011001101;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101011001100000011001011;
#10000;
	data_in <= 24'b101011001100000011001011;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101011011100001011001011;
#10000;
	data_in <= 24'b101010001011111011001000;
#10000;
	data_in <= 24'b101001111011110111001000;
#10000;
	data_in <= 24'b101001111011110111001000;
#10000;
	data_in <= 24'b101001111011110111000111;
#10000;
	data_in <= 24'b101001111011110111000111;
#10000;
	data_in <= 24'b101001111011110111001000;
#10000;
	data_in <= 24'b101001111011110111000111;
#10000;
	data_in <= 24'b101010001011111011001000;
#10000;
	data_in <= 24'b101001011011101111000101;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b101001001011101011000100;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
	data_in <= 24'b101000111011100111000100;
#10000;
	data_in <= 24'b101000101011100111000100;
#10000;
	data_in <= 24'b101000101011100111000100;
#10000;
	data_in <= 24'b101000101011100111000100;
#10000;
	data_in <= 24'b101000111011100111000100;
#10000;
	data_in <= 24'b101000111011100111000100;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101001001011101111000101;
#10000;
	data_in <= 24'b101000111011101111000101;
#10000;
	data_in <= 24'b101000111011101111000101;
#10000;
	data_in <= 24'b101000111011101111000101;
#10000;
	data_in <= 24'b101000111011101111000101;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
	data_in <= 24'b101001001011101111000101;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101101101100101111010101;
#10000;
	data_in <= 24'b101101011100101011010101;
#10000;
	data_in <= 24'b101100101100011011001111;
#10000;
	data_in <= 24'b101010101011010110110101;
#10000;
	data_in <= 24'b101000001001100110001000;
#10000;
	data_in <= 24'b100111101000100001101000;
#10000;
	data_in <= 24'b101001001000101001100110;
#10000;
	data_in <= 24'b101010101001001001101101;
#10000;
	data_in <= 24'b101100101100010011001110;
#10000;
	data_in <= 24'b101100101100010111001110;
#10000;
	data_in <= 24'b101100101100011011001111;
#10000;
	data_in <= 24'b101100111100100011010011;
#10000;
	data_in <= 24'b101100001100011011010010;
#10000;
	data_in <= 24'b101001111011000110110000;
#10000;
	data_in <= 24'b100111011001000001110111;
#10000;
	data_in <= 24'b100000000111001101011011;
#10000;
	data_in <= 24'b101011101100001011001100;
#10000;
	data_in <= 24'b101011111100001111001100;
#10000;
	data_in <= 24'b101011111100001111001101;
#10000;
	data_in <= 24'b101011111100001111001100;
#10000;
	data_in <= 24'b101011111100001111001100;
#10000;
	data_in <= 24'b101100001100011011010010;
#10000;
	data_in <= 24'b101011001011111011000100;
#10000;
	data_in <= 24'b010111000110110001110100;
#10000;
	data_in <= 24'b101010011011111111001001;
#10000;
	data_in <= 24'b101010101100000011001010;
#10000;
	data_in <= 24'b101011001100000111001010;
#10000;
	data_in <= 24'b101011011100000111001100;
#10000;
	data_in <= 24'b101011101100001011001011;
#10000;
	data_in <= 24'b101011001100000011001000;
#10000;
	data_in <= 24'b101011011100001011001101;
#10000;
	data_in <= 24'b101010011011111011001000;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101001111011110011000111;
#10000;
	data_in <= 24'b101010001011110111001000;
#10000;
	data_in <= 24'b101010101011111111001001;
#10000;
	data_in <= 24'b101010111100000011001010;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101010101011111011000111;
#10000;
	data_in <= 24'b101011011100000111001010;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101001101011110011000111;
#10000;
	data_in <= 24'b101001111011110111000111;
#10000;
	data_in <= 24'b101010011011111011001001;
#10000;
	data_in <= 24'b101010111100000011001001;
#10000;
	data_in <= 24'b101010111100000011001010;
#10000;
	data_in <= 24'b101001111011110011000110;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
	data_in <= 24'b101000001011100011000100;
#10000;
	data_in <= 24'b101000001011100011000011;
#10000;
	data_in <= 24'b101000011011100111000100;
#10000;
	data_in <= 24'b101000101011100111000100;
#10000;
	data_in <= 24'b101000101011101011000101;
#10000;
	data_in <= 24'b101001111011110111001000;
#10000;
	data_in <= 24'b101010101011111111001000;
#10000;
	data_in <= 24'b101000001011100011000011;
#10000;
	data_in <= 24'b101011111100000111001010;
#10000;
	data_in <= 24'b110001111101001011010111;
#10000;
	data_in <= 24'b110100111101101111011111;
#10000;
	data_in <= 24'b110100011101101011011110;
#10000;
	data_in <= 24'b110000101100111111010101;
#10000;
	data_in <= 24'b101010101011111111001000;
#10000;
	data_in <= 24'b101001001011101111000110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000111000110001101000;
#10000;
	data_in <= 24'b100110001000010101100101;
#10000;
	data_in <= 24'b100110011000010101100101;
#10000;
	data_in <= 24'b101000111000101101100110;
#10000;
	data_in <= 24'b101001111000110101100111;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101000111000100101100100;
#10000;
	data_in <= 24'b010110110110000001011110;
#10000;
	data_in <= 24'b010100000101110001100001;
#10000;
	data_in <= 24'b010101010101111101100010;
#10000;
	data_in <= 24'b011001010110100001100010;
#10000;
	data_in <= 24'b100001110111101101100011;
#10000;
	data_in <= 24'b101001011000110101100111;
#10000;
	data_in <= 24'b101001101000111001101000;
#10000;
	data_in <= 24'b101001011000110101101000;
#10000;
	data_in <= 24'b001000110011101001001010;
#10000;
	data_in <= 24'b001111000101000101011111;
#10000;
	data_in <= 24'b001111110101010001100011;
#10000;
	data_in <= 24'b001111000101001001100001;
#10000;
	data_in <= 24'b001111100101000001011011;
#10000;
	data_in <= 24'b011001110110011001011101;
#10000;
	data_in <= 24'b101000101000101101101001;
#10000;
	data_in <= 24'b101010001001000001101010;
#10000;
	data_in <= 24'b010110010110110001111000;
#10000;
	data_in <= 24'b001010010011111101001100;
#10000;
	data_in <= 24'b001110110101000001011101;
#10000;
	data_in <= 24'b001111000101000101011101;
#10000;
	data_in <= 24'b001101110100110001011001;
#10000;
	data_in <= 24'b001010110100000101010001;
#10000;
	data_in <= 24'b010110000101101101010110;
#10000;
	data_in <= 24'b101001011000110101101011;
#10000;
	data_in <= 24'b101001111011101111000101;
#10000;
	data_in <= 24'b010001010101101101101000;
#10000;
	data_in <= 24'b000111110011011001000101;
#10000;
	data_in <= 24'b001011110100011001010100;
#10000;
	data_in <= 24'b001011100100010101010010;
#10000;
	data_in <= 24'b001011000100001001001111;
#10000;
	data_in <= 24'b000111100011010101000101;
#10000;
	data_in <= 24'b011000100110000101010110;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b100101001010100110110100;
#10000;
	data_in <= 24'b001001000011101101001000;
#10000;
	data_in <= 24'b000110000011000100111111;
#10000;
	data_in <= 24'b001000100011101001001000;
#10000;
	data_in <= 24'b001000110011101001001000;
#10000;
	data_in <= 24'b000111100011010001000011;
#10000;
	data_in <= 24'b000111000010111100111100;
#10000;
	data_in <= 24'b101001011011101011000011;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b011010011000000010001011;
#10000;
	data_in <= 24'b000001100001111000101110;
#10000;
	data_in <= 24'b000101010010111000111101;
#10000;
	data_in <= 24'b000110000011000000111111;
#10000;
	data_in <= 24'b000110010011000000111110;
#10000;
	data_in <= 24'b000010110010001100110011;
#10000;
	data_in <= 24'b101001111011110011000110;
#10000;
	data_in <= 24'b101001011011101011000100;
#10000;
	data_in <= 24'b100111111011010010111111;
#10000;
	data_in <= 24'b001010010100000001001110;
#10000;
	data_in <= 24'b000000100001100100101000;
#10000;
	data_in <= 24'b000100000010101000111001;
#10000;
	data_in <= 24'b000011110010100000110111;
#10000;
	data_in <= 24'b000010010010000100110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000101000100001100011;
#10000;
	data_in <= 24'b101000011000011101100001;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b100111111000010001011111;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b100111011000000101011101;
#10000;
	data_in <= 24'b100110111000000001011010;
#10000;
	data_in <= 24'b100110010111111101011000;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
	data_in <= 24'b101001011000101101100110;
#10000;
	data_in <= 24'b101001001000101101100100;
#10000;
	data_in <= 24'b101000101000100101100010;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b100111111000010101011111;
#10000;
	data_in <= 24'b100111101000001101011101;
#10000;
	data_in <= 24'b100111001000001001011011;
#10000;
	data_in <= 24'b101001111000111101101001;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101001101000111001101000;
#10000;
	data_in <= 24'b101001011000110101100110;
#10000;
	data_in <= 24'b101000111000101001100100;
#10000;
	data_in <= 24'b101000101000100001100011;
#10000;
	data_in <= 24'b101000001000011101100000;
#10000;
	data_in <= 24'b100111111000010101011110;
#10000;
	data_in <= 24'b101010101001001001101101;
#10000;
	data_in <= 24'b101010011001000101101100;
#10000;
	data_in <= 24'b101010001001000001101010;
#10000;
	data_in <= 24'b101001111000111101101000;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101001001000101101100101;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b101000101000100001100001;
#10000;
	data_in <= 24'b101011101001010001110000;
#10000;
	data_in <= 24'b101010111001001101101111;
#10000;
	data_in <= 24'b101010111001001101101110;
#10000;
	data_in <= 24'b101010011001001001101100;
#10000;
	data_in <= 24'b101010001001000101101010;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101001101000110001100111;
#10000;
	data_in <= 24'b101001001000101001100100;
#10000;
	data_in <= 24'b100001100111100101100001;
#10000;
	data_in <= 24'b101100101001100101110011;
#10000;
	data_in <= 24'b101011011001010101110001;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b101010111001010001101110;
#10000;
	data_in <= 24'b101010011001000001101011;
#10000;
	data_in <= 24'b101010001000111001101010;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b001111010100010001000100;
#10000;
	data_in <= 24'b101011111001011101110011;
#10000;
	data_in <= 24'b101011111001100001110010;
#10000;
	data_in <= 24'b101011111001011101110001;
#10000;
	data_in <= 24'b101011101001011001110000;
#10000;
	data_in <= 24'b101011001001010001101110;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101010011001000001101001;
#10000;
	data_in <= 24'b000011000010000000101100;
#10000;
	data_in <= 24'b100010100111110001100100;
#10000;
	data_in <= 24'b101110011001111101111001;
#10000;
	data_in <= 24'b101100001001100001110100;
#10000;
	data_in <= 24'b101100011001100001110010;
#10000;
	data_in <= 24'b101011111001011001110001;
#10000;
	data_in <= 24'b101011101001010001101111;
#10000;
	data_in <= 24'b101011001001001001101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100101110111110101010110;
#10000;
	data_in <= 24'b100101100111101101010011;
#10000;
	data_in <= 24'b100101000111100101010001;
#10000;
	data_in <= 24'b100100100111011101001111;
#10000;
	data_in <= 24'b100100010111010101001101;
#10000;
	data_in <= 24'b100011100111001101001100;
#10000;
	data_in <= 24'b100011000111000001001000;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100110101000000001011010;
#10000;
	data_in <= 24'b100110010111111001010111;
#10000;
	data_in <= 24'b100101110111110101010100;
#10000;
	data_in <= 24'b100101010111101001010011;
#10000;
	data_in <= 24'b100100110111100001010000;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b100011110111010001001011;
#10000;
	data_in <= 24'b100011010111001001001000;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100110100111111101011000;
#10000;
	data_in <= 24'b100110000111110101010110;
#10000;
	data_in <= 24'b100101010111101101010100;
#10000;
	data_in <= 24'b100100110111100101010001;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b100100000111010001001100;
#10000;
	data_in <= 24'b101000001000011001011111;
#10000;
	data_in <= 24'b100111101000010001011101;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100110100111111101011000;
#10000;
	data_in <= 24'b100101110111110101010110;
#10000;
	data_in <= 24'b100101010111101101010011;
#10000;
	data_in <= 24'b100100110111100101010000;
#10000;
	data_in <= 24'b100100010111011001001110;
#10000;
	data_in <= 24'b101000111000100101100010;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b100111101000001101011101;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100110101000000001011001;
#10000;
	data_in <= 24'b100110000111111001010110;
#10000;
	data_in <= 24'b100101010111101101010011;
#10000;
	data_in <= 24'b100100110111100001010001;
#10000;
	data_in <= 24'b101001011000110001100101;
#10000;
	data_in <= 24'b101000111000101001100011;
#10000;
	data_in <= 24'b101000011000011101100000;
#10000;
	data_in <= 24'b100111011000010001011101;
#10000;
	data_in <= 24'b100111001000001001011011;
#10000;
	data_in <= 24'b100110101000000001011001;
#10000;
	data_in <= 24'b100110000111111001010110;
#10000;
	data_in <= 24'b100101010111101001010011;
#10000;
	data_in <= 24'b101001111000111001100111;
#10000;
	data_in <= 24'b101001101000110101100101;
#10000;
	data_in <= 24'b101000111000101001100010;
#10000;
	data_in <= 24'b101000001000011101100000;
#10000;
	data_in <= 24'b100111101000010101011101;
#10000;
	data_in <= 24'b100111001000001101011011;
#10000;
	data_in <= 24'b100110101000000001011000;
#10000;
	data_in <= 24'b100110000111110101010110;
#10000;
	data_in <= 24'b101010101001000001101011;
#10000;
	data_in <= 24'b101010001000111001100111;
#10000;
	data_in <= 24'b101001111000110001100110;
#10000;
	data_in <= 24'b101001001000100101100011;
#10000;
	data_in <= 24'b101000011000011101100001;
#10000;
	data_in <= 24'b100111101000010001011101;
#10000;
	data_in <= 24'b100111011000000101011011;
#10000;
	data_in <= 24'b100110100111111001011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010010110110001000100;
#10000;
	data_in <= 24'b100001110110101001000001;
#10000;
	data_in <= 24'b100001010110011100111110;
#10000;
	data_in <= 24'b100000100110010100111100;
#10000;
	data_in <= 24'b011111110110001000111001;
#10000;
	data_in <= 24'b011111010101111100110110;
#10000;
	data_in <= 24'b011110110101110100110011;
#10000;
	data_in <= 24'b011110000101101000110001;
#10000;
	data_in <= 24'b100010110110111101000110;
#10000;
	data_in <= 24'b100010010110110001000011;
#10000;
	data_in <= 24'b100001110110101001000001;
#10000;
	data_in <= 24'b100001000110011100111110;
#10000;
	data_in <= 24'b100000010110010100111011;
#10000;
	data_in <= 24'b011111110110001000111000;
#10000;
	data_in <= 24'b011111010101111100110101;
#10000;
	data_in <= 24'b011110100101110100110010;
#10000;
	data_in <= 24'b100011100111001001001001;
#10000;
	data_in <= 24'b100010110110111001000101;
#10000;
	data_in <= 24'b100010010110110001000011;
#10000;
	data_in <= 24'b100001110110101001000001;
#10000;
	data_in <= 24'b100000110110011100111110;
#10000;
	data_in <= 24'b100000000110010000111010;
#10000;
	data_in <= 24'b011111100110000100110111;
#10000;
	data_in <= 24'b011111000110000000110100;
#10000;
	data_in <= 24'b100011110111010001001011;
#10000;
	data_in <= 24'b100011010111000101001000;
#10000;
	data_in <= 24'b100010110110111001000101;
#10000;
	data_in <= 24'b100010000110101101000010;
#10000;
	data_in <= 24'b100001100110100101000000;
#10000;
	data_in <= 24'b100000110110011100111100;
#10000;
	data_in <= 24'b100000000110001100111001;
#10000;
	data_in <= 24'b011111010110000000110101;
#10000;
	data_in <= 24'b100100010111010101001101;
#10000;
	data_in <= 24'b100011110111001101001011;
#10000;
	data_in <= 24'b100011010111000001000111;
#10000;
	data_in <= 24'b100010100110110101000101;
#10000;
	data_in <= 24'b100001110110101101000010;
#10000;
	data_in <= 24'b100001000110100000111111;
#10000;
	data_in <= 24'b100000010110010000111011;
#10000;
	data_in <= 24'b011111100110000100111000;
#10000;
	data_in <= 24'b100100110111100001001111;
#10000;
	data_in <= 24'b100100010111011001001101;
#10000;
	data_in <= 24'b100011110111001101001010;
#10000;
	data_in <= 24'b100011000111000001000111;
#10000;
	data_in <= 24'b100010000110110101000011;
#10000;
	data_in <= 24'b100001010110101001000000;
#10000;
	data_in <= 24'b100000100110011000111101;
#10000;
	data_in <= 24'b011111110110001100111001;
#10000;
	data_in <= 24'b100101010111101001010010;
#10000;
	data_in <= 24'b100100110111011101001111;
#10000;
	data_in <= 24'b100100000111010101001100;
#10000;
	data_in <= 24'b100011110111001001001001;
#10000;
	data_in <= 24'b100010110110111001000101;
#10000;
	data_in <= 24'b100001110110110001000001;
#10000;
	data_in <= 24'b100001000110100000111110;
#10000;
	data_in <= 24'b100000010110010000111011;
#10000;
	data_in <= 24'b100110000111110001010100;
#10000;
	data_in <= 24'b100101010111100101010001;
#10000;
	data_in <= 24'b100100110111011001001110;
#10000;
	data_in <= 24'b100100010111010001001011;
#10000;
	data_in <= 24'b100011010111000001000111;
#10000;
	data_in <= 24'b100010010110110101000011;
#10000;
	data_in <= 24'b100001110110101001000000;
#10000;
	data_in <= 24'b100001000110011000111101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100001000110011100111110;
#10000;
	data_in <= 24'b100001110110101101000010;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100011110111001001001001;
#10000;
	data_in <= 24'b100100100111010101001100;
#10000;
	data_in <= 24'b100101010111100001010000;
#10000;
	data_in <= 24'b100101110111101101010011;
#10000;
	data_in <= 24'b100110100111111001010110;
#10000;
	data_in <= 24'b100001100110100101000000;
#10000;
	data_in <= 24'b100010000110110101000100;
#10000;
	data_in <= 24'b100011000111000001001000;
#10000;
	data_in <= 24'b100100010111010001001011;
#10000;
	data_in <= 24'b100100110111011101001110;
#10000;
	data_in <= 24'b100101100111101001010010;
#10000;
	data_in <= 24'b100110000111110101010101;
#10000;
	data_in <= 24'b100110110111111101011000;
#10000;
	data_in <= 24'b100001110110101001000010;
#10000;
	data_in <= 24'b100010010110111001000101;
#10000;
	data_in <= 24'b100011100111001001001001;
#10000;
	data_in <= 24'b100100100111010101001101;
#10000;
	data_in <= 24'b100101000111100101001111;
#10000;
	data_in <= 24'b100101110111110001010011;
#10000;
	data_in <= 24'b100110100111111101010111;
#10000;
	data_in <= 24'b100111001000001001011010;
#10000;
	data_in <= 24'b100001110110101101000011;
#10000;
	data_in <= 24'b100010100110111101000111;
#10000;
	data_in <= 24'b100011110111001101001011;
#10000;
	data_in <= 24'b100100110111011001001110;
#10000;
	data_in <= 24'b100101100111101001010010;
#10000;
	data_in <= 24'b100110010111111001010110;
#10000;
	data_in <= 24'b100110111000000001011001;
#10000;
	data_in <= 24'b100111101000001101011100;
#10000;
	data_in <= 24'b100010000110110101000101;
#10000;
	data_in <= 24'b100010110111000101001001;
#10000;
	data_in <= 24'b100100000111010001001101;
#10000;
	data_in <= 24'b100101000111011101010000;
#10000;
	data_in <= 24'b100101110111110001010100;
#10000;
	data_in <= 24'b100110100111111101011000;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100111111000010001011111;
#10000;
	data_in <= 24'b100010010110111001000110;
#10000;
	data_in <= 24'b100011010111001101001010;
#10000;
	data_in <= 24'b100100100111011101001110;
#10000;
	data_in <= 24'b100101010111101001010001;
#10000;
	data_in <= 24'b100110000111110101010101;
#10000;
	data_in <= 24'b100110111000000101011001;
#10000;
	data_in <= 24'b100111101000010001011100;
#10000;
	data_in <= 24'b101000011000011101100000;
#10000;
	data_in <= 24'b100010100111000001001000;
#10000;
	data_in <= 24'b100011100111010101001100;
#10000;
	data_in <= 24'b100100110111100001001111;
#10000;
	data_in <= 24'b100101100111101101010011;
#10000;
	data_in <= 24'b100110010111111001010110;
#10000;
	data_in <= 24'b100111011000001001011011;
#10000;
	data_in <= 24'b100111111000010101011110;
#10000;
	data_in <= 24'b101000101000100001100010;
#10000;
	data_in <= 24'b100010110111000001001001;
#10000;
	data_in <= 24'b100011110111010101001101;
#10000;
	data_in <= 24'b100101000111100101010000;
#10000;
	data_in <= 24'b100110000111101101010100;
#10000;
	data_in <= 24'b100110101000000001011000;
#10000;
	data_in <= 24'b100111101000001101011100;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100111001000000001011001;
#10000;
	data_in <= 24'b100111101000010001011100;
#10000;
	data_in <= 24'b101000011000011101011111;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b101001011000101101100101;
#10000;
	data_in <= 24'b101010001000111001100111;
#10000;
	data_in <= 24'b101010101001000001101001;
#10000;
	data_in <= 24'b101011011001001101101101;
#10000;
	data_in <= 24'b100111011000001101011100;
#10000;
	data_in <= 24'b101000001000011101011111;
#10000;
	data_in <= 24'b101000101000100101100010;
#10000;
	data_in <= 24'b101001001000101101100101;
#10000;
	data_in <= 24'b101001111000110101101000;
#10000;
	data_in <= 24'b101010101001000001101010;
#10000;
	data_in <= 24'b101011011001010001101101;
#10000;
	data_in <= 24'b101011101001010101101111;
#10000;
	data_in <= 24'b100111111000010101011101;
#10000;
	data_in <= 24'b101000101000100101100001;
#10000;
	data_in <= 24'b101001001000101101100100;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101010011000111101101011;
#10000;
	data_in <= 24'b101011001001001001101101;
#10000;
	data_in <= 24'b101011101001010101101111;
#10000;
	data_in <= 24'b101100001001011101110001;
#10000;
	data_in <= 24'b101000001000011001011111;
#10000;
	data_in <= 24'b101000111000101001100011;
#10000;
	data_in <= 24'b101001011000110001100110;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101010111001000101101100;
#10000;
	data_in <= 24'b101011101001010001101111;
#10000;
	data_in <= 24'b101100001001011101110001;
#10000;
	data_in <= 24'b101100101001100101110100;
#10000;
	data_in <= 24'b101000101000100001100010;
#10000;
	data_in <= 24'b101001011000101101100110;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101010011001000001101011;
#10000;
	data_in <= 24'b101011011001001101101110;
#10000;
	data_in <= 24'b101011111001011001110001;
#10000;
	data_in <= 24'b101100101001100001110011;
#10000;
	data_in <= 24'b101101001001101101110110;
#10000;
	data_in <= 24'b101000111000100101100100;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101011001001001101101100;
#10000;
	data_in <= 24'b101011101001010101110000;
#10000;
	data_in <= 24'b101100001001100001110010;
#10000;
	data_in <= 24'b101100111001101101110101;
#10000;
	data_in <= 24'b101101101001110101111000;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101001111000111101101000;
#10000;
	data_in <= 24'b101010101001001001101100;
#10000;
	data_in <= 24'b101011011001010101101111;
#10000;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b101100101001101001110100;
#10000;
	data_in <= 24'b101101011001110101110111;
#10000;
	data_in <= 24'b101101111001111101111011;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101010111001001101101101;
#10000;
	data_in <= 24'b101011101001011001110001;
#10000;
	data_in <= 24'b101100011001100001110100;
#10000;
	data_in <= 24'b101101001001101101110110;
#10000;
	data_in <= 24'b101101111001111001111001;
#10000;
	data_in <= 24'b101110001010000001111100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101011101001010001101111;
#10000;
	data_in <= 24'b101100001001011001110001;
#10000;
	data_in <= 24'b101100011001100001110011;
#10000;
	data_in <= 24'b101100101001101001110101;
#10000;
	data_in <= 24'b101101001001110001110111;
#10000;
	data_in <= 24'b101101011001111001111000;
#10000;
	data_in <= 24'b101101111001111101111011;
#10000;
	data_in <= 24'b101110001010000101111101;
#10000;
	data_in <= 24'b101100001001011101110001;
#10000;
	data_in <= 24'b101100101001100101110011;
#10000;
	data_in <= 24'b101100111001101101110110;
#10000;
	data_in <= 24'b101101011001110101111001;
#10000;
	data_in <= 24'b101101101001111101111010;
#10000;
	data_in <= 24'b101101111010000101111100;
#10000;
	data_in <= 24'b101110011010001001111110;
#10000;
	data_in <= 24'b101110111010001101111111;
#10000;
	data_in <= 24'b101100101001100101110100;
#10000;
	data_in <= 24'b101101001001110001110110;
#10000;
	data_in <= 24'b101101011001110101111001;
#10000;
	data_in <= 24'b101101111010000001111011;
#10000;
	data_in <= 24'b101110001010000101111100;
#10000;
	data_in <= 24'b101110101010001101111110;
#10000;
	data_in <= 24'b101110111010010010000001;
#10000;
	data_in <= 24'b101111101010011010000010;
#10000;
	data_in <= 24'b101101001001101101110111;
#10000;
	data_in <= 24'b101101101001111001111000;
#10000;
	data_in <= 24'b101101111001111101111011;
#10000;
	data_in <= 24'b101110011010000101111101;
#10000;
	data_in <= 24'b101110111010001101111110;
#10000;
	data_in <= 24'b101110111010010010000000;
#10000;
	data_in <= 24'b101111011010011010000011;
#10000;
	data_in <= 24'b110000001010100010000101;
#10000;
	data_in <= 24'b101101101001110101111001;
#10000;
	data_in <= 24'b101101111001111101111010;
#10000;
	data_in <= 24'b101110011010000101111110;
#10000;
	data_in <= 24'b101110111010001110000000;
#10000;
	data_in <= 24'b101111001010010110000001;
#10000;
	data_in <= 24'b101111011010011010000011;
#10000;
	data_in <= 24'b110000001010100010000101;
#10000;
	data_in <= 24'b110000101010101010000111;
#10000;
	data_in <= 24'b101101111001111101111010;
#10000;
	data_in <= 24'b101110011010000101111101;
#10000;
	data_in <= 24'b101110111010001110000000;
#10000;
	data_in <= 24'b101111001010011010000001;
#10000;
	data_in <= 24'b101111101010100010000011;
#10000;
	data_in <= 24'b101111111010100110000101;
#10000;
	data_in <= 24'b110000101010101110000111;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b101110011010000101111100;
#10000;
	data_in <= 24'b101110111010001101111110;
#10000;
	data_in <= 24'b101111001010010110000001;
#10000;
	data_in <= 24'b101111101010100010000100;
#10000;
	data_in <= 24'b110000001010101010000110;
#10000;
	data_in <= 24'b110000011010101110000111;
#10000;
	data_in <= 24'b110001001010110010001010;
#10000;
	data_in <= 24'b110001101010111010001100;
#10000;
	data_in <= 24'b101110101010001001111110;
#10000;
	data_in <= 24'b101111001010010110000000;
#10000;
	data_in <= 24'b101111101010011110000011;
#10000;
	data_in <= 24'b110000001010100110000110;
#10000;
	data_in <= 24'b110000011010101110000111;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110001011010111010001011;
#10000;
	data_in <= 24'b110001111010111110001101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101110101010001001111110;
#10000;
	data_in <= 24'b101110111010001101111111;
#10000;
	data_in <= 24'b101111001010010010000000;
#10000;
	data_in <= 24'b101111011010010110000010;
#10000;
	data_in <= 24'b101111101010011010000011;
#10000;
	data_in <= 24'b101101011001111101111111;
#10000;
	data_in <= 24'b001010010011001000110111;
#10000;
	data_in <= 24'b000000000001001000100011;
#10000;
	data_in <= 24'b101111001010010010000000;
#10000;
	data_in <= 24'b101111101010011010000010;
#10000;
	data_in <= 24'b101111101010011110000011;
#10000;
	data_in <= 24'b101111111010100010000100;
#10000;
	data_in <= 24'b110000111010101110000111;
#10000;
	data_in <= 24'b101000101001001001110111;
#10000;
	data_in <= 24'b000011000001110000101000;
#10000;
	data_in <= 24'b000000000001010000100100;
#10000;
	data_in <= 24'b101111111010011110000011;
#10000;
	data_in <= 24'b110000001010100110000101;
#10000;
	data_in <= 24'b110000011010101010000110;
#10000;
	data_in <= 24'b110000011010101010000111;
#10000;
	data_in <= 24'b110001111010111110001011;
#10000;
	data_in <= 24'b100100111000011001101111;
#10000;
	data_in <= 24'b000000100001001000100010;
#10000;
	data_in <= 24'b000000000001010000100101;
#10000;
	data_in <= 24'b110000011010100110000110;
#10000;
	data_in <= 24'b110000101010101010000111;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110010101011001010001110;
#10000;
	data_in <= 24'b100100001000001101101111;
#10000;
	data_in <= 24'b000000010001000000100000;
#10000;
	data_in <= 24'b000000000001001000100011;
#10000;
	data_in <= 24'b110000111010101110001000;
#10000;
	data_in <= 24'b110001001010110010001001;
#10000;
	data_in <= 24'b110001011010111010001100;
#10000;
	data_in <= 24'b110001001010111010001100;
#10000;
	data_in <= 24'b110010111011001110010000;
#10000;
	data_in <= 24'b100110001000101001110011;
#10000;
	data_in <= 24'b000000110000111100011110;
#10000;
	data_in <= 24'b000000000000111100100000;
#10000;
	data_in <= 24'b110001011010110110001010;
#10000;
	data_in <= 24'b110001101010111110001011;
#10000;
	data_in <= 24'b110001101011000010001110;
#10000;
	data_in <= 24'b110001111011000110001110;
#10000;
	data_in <= 24'b110010111011010010010001;
#10000;
	data_in <= 24'b101011001001101110000000;
#10000;
	data_in <= 24'b000011110001011000100010;
#10000;
	data_in <= 24'b000000000000100100011011;
#10000;
	data_in <= 24'b110001101010111110001100;
#10000;
	data_in <= 24'b110001111011000010001110;
#10000;
	data_in <= 24'b110010001011001010010000;
#10000;
	data_in <= 24'b110010011011001110010010;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110000111011000010010001;
#10000;
	data_in <= 24'b001100100011000000110101;
#10000;
	data_in <= 24'b000000010000000100010100;
#10000;
	data_in <= 24'b110010011011000110001110;
#10000;
	data_in <= 24'b110010101011001010010000;
#10000;
	data_in <= 24'b110010101011010010010010;
#10000;
	data_in <= 24'b110010111011010110010011;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110100011011110010011001;
#10000;
	data_in <= 24'b011110010110111001100010;
#10000;
	data_in <= 24'b000000000000000000001110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001100001111100101110;
#10000;
	data_in <= 24'b000010000010001000110010;
#10000;
	data_in <= 24'b000000010001010100100100;
#10000;
	data_in <= 24'b001100000100011001010011;
#10000;
	data_in <= 24'b101000101011011111000010;
#10000;
	data_in <= 24'b101000111011100111000011;
#10000;
	data_in <= 24'b101001111011110011000111;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b000000010001100100101001;
#10000;
	data_in <= 24'b000000100001101100101011;
#10000;
	data_in <= 24'b000000000001001000100010;
#10000;
	data_in <= 24'b011010000111111010001011;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101000111011100111000011;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b110001001100111111010100;
#10000;
	data_in <= 24'b000000100001100100101001;
#10000;
	data_in <= 24'b000000000001001000100010;
#10000;
	data_in <= 24'b000101100010100100111001;
#10000;
	data_in <= 24'b100011011010001110101110;
#10000;
	data_in <= 24'b101001011011101011000100;
#10000;
	data_in <= 24'b101000101011100011000011;
#10000;
	data_in <= 24'b101011101100000111001010;
#10000;
	data_in <= 24'b111010001110100011101000;
#10000;
	data_in <= 24'b000000110001011100101000;
#10000;
	data_in <= 24'b000000000000101100011100;
#10000;
	data_in <= 24'b001101110100101101011001;
#10000;
	data_in <= 24'b100111101011010110111111;
#10000;
	data_in <= 24'b101000101011011111000001;
#10000;
	data_in <= 24'b101000011011100011000010;
#10000;
	data_in <= 24'b110000101100111011010011;
#10000;
	data_in <= 24'b111100011111000011101111;
#10000;
	data_in <= 24'b000000010001001100100100;
#10000;
	data_in <= 24'b000000000000101000011011;
#10000;
	data_in <= 24'b010101100110101001110111;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101000011011011011000000;
#10000;
	data_in <= 24'b101000011011100011000011;
#10000;
	data_in <= 24'b110011001101010111011001;
#10000;
	data_in <= 24'b111100011111000111110000;
#10000;
	data_in <= 24'b000000000000110000011100;
#10000;
	data_in <= 24'b000001000000111000011111;
#10000;
	data_in <= 24'b011011111000010010010000;
#10000;
	data_in <= 24'b101001111011110111000111;
#10000;
	data_in <= 24'b101000101011011111000001;
#10000;
	data_in <= 24'b101000101011100111000011;
#10000;
	data_in <= 24'b110010111101010011011000;
#10000;
	data_in <= 24'b111100001110111111101111;
#10000;
	data_in <= 24'b000000000000010000010111;
#10000;
	data_in <= 24'b000011100001001000100100;
#10000;
	data_in <= 24'b100000011001011010100011;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101001001011100011000011;
#10000;
	data_in <= 24'b101000101011101011000101;
#10000;
	data_in <= 24'b110001001100111111010101;
#10000;
	data_in <= 24'b111100001110111111101111;
#10000;
	data_in <= 24'b000000100000001000010000;
#10000;
	data_in <= 24'b000101100001101000101100;
#10000;
	data_in <= 24'b100011001010001010101110;
#10000;
	data_in <= 24'b101001001011101011000100;
#10000;
	data_in <= 24'b101001011011101011000011;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101110011100100011001111;
#10000;
	data_in <= 24'b111011101110110111101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001011101000011010101;
#10000;
	data_in <= 24'b111010111110101111101011;
#10000;
	data_in <= 24'b111101111111011011110100;
#10000;
	data_in <= 24'b111110101111100111111000;
#10000;
	data_in <= 24'b111111001111101111111010;
#10000;
	data_in <= 24'b111111001111101011111010;
#10000;
	data_in <= 24'b111010111110111011101111;
#10000;
	data_in <= 24'b101110101100100111010001;
#10000;
	data_in <= 24'b111100101111000011110000;
#10000;
	data_in <= 24'b111101001111010011110011;
#10000;
	data_in <= 24'b111100111111001111110011;
#10000;
	data_in <= 24'b111100111111010011110100;
#10000;
	data_in <= 24'b111100111111010011110100;
#10000;
	data_in <= 24'b111101111111011111111000;
#10000;
	data_in <= 24'b111111111111111111111110;
#10000;
	data_in <= 24'b111101101111011011110110;
#10000;
	data_in <= 24'b111100111111001011110010;
#10000;
	data_in <= 24'b111100011111000111110001;
#10000;
	data_in <= 24'b111100101111001011110010;
#10000;
	data_in <= 24'b111110011111100111111001;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111110101111101011111010;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111100001111000011110000;
#10000;
	data_in <= 24'b111100011111000111110001;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b110100011101001011010101;
#10000;
	data_in <= 24'b011110111000000010000110;
#10000;
	data_in <= 24'b101111111100000111000100;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111111001111110011111100;
#10000;
	data_in <= 24'b111100101111001011110010;
#10000;
	data_in <= 24'b111010101110101111101011;
#10000;
	data_in <= 24'b101100111011010110110111;
#10000;
	data_in <= 24'b100011001001000010010101;
#10000;
	data_in <= 24'b000001110001000100011011;
#10000;
	data_in <= 24'b000101100001111000101000;
#10000;
	data_in <= 24'b101011001010111010110001;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111101111111011111110111;
#10000;
	data_in <= 24'b110100111101010011010101;
#10000;
	data_in <= 24'b001100000011010100111010;
#10000;
	data_in <= 24'b000101010010000000100111;
#10000;
	data_in <= 24'b000100000001110000100011;
#10000;
	data_in <= 24'b000000000000001100001001;
#10000;
	data_in <= 24'b010111000101111001100001;
#10000;
	data_in <= 24'b111000001110001111100101;
#10000;
	data_in <= 24'b111110001111100011110111;
#10000;
	data_in <= 24'b110111111101111011011101;
#10000;
	data_in <= 24'b001010110010111000110001;
#10000;
	data_in <= 24'b000111000010010000101001;
#10000;
	data_in <= 24'b001110110100010101001011;
#10000;
	data_in <= 24'b010010100101001101011001;
#10000;
	data_in <= 24'b010110010110001101101001;
#10000;
	data_in <= 24'b010001010101110101101000;
#10000;
	data_in <= 24'b111001101110100111101011;
#10000;
	data_in <= 24'b110101101101110111100010;
#10000;
	data_in <= 24'b101010101011011010111101;
#10000;
	data_in <= 24'b101100111100000111001001;
#10000;
	data_in <= 24'b110010011101011111011111;
#10000;
	data_in <= 24'b101110001100100111010010;
#10000;
	data_in <= 24'b001110100101010001100001;
#10000;
	data_in <= 24'b000111010011101001001000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000011011100111000100;
#10000;
	data_in <= 24'b101001011011110011000110;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101001011011101111000110;
#10000;
	data_in <= 24'b101001001011101111000110;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b101101101100011111001111;
#10000;
	data_in <= 24'b101000101011100111000100;
#10000;
	data_in <= 24'b101001101011110011000111;
#10000;
	data_in <= 24'b101001011011110011000110;
#10000;
	data_in <= 24'b101001011011110011000110;
#10000;
	data_in <= 24'b101001101011110011000111;
#10000;
	data_in <= 24'b101000101011101011000101;
#10000;
	data_in <= 24'b110001111101000111010110;
#10000;
	data_in <= 24'b111000111110100011101011;
#10000;
	data_in <= 24'b101001001011101011000101;
#10000;
	data_in <= 24'b101001101011101111000110;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101000111011101011000101;
#10000;
	data_in <= 24'b101100011100001011001010;
#10000;
	data_in <= 24'b111010101110101011101010;
#10000;
	data_in <= 24'b111101101111011111110111;
#10000;
	data_in <= 24'b101110011100101011010010;
#10000;
	data_in <= 24'b101010001011111111001010;
#10000;
	data_in <= 24'b101011101100010011001101;
#10000;
	data_in <= 24'b101011011100001111001101;
#10000;
	data_in <= 24'b101010001011111111001010;
#10000;
	data_in <= 24'b110001101101000011010101;
#10000;
	data_in <= 24'b111011111110111011101101;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b101110011100100011001111;
#10000;
	data_in <= 24'b100100001010100010110011;
#10000;
	data_in <= 24'b100011011010001110101101;
#10000;
	data_in <= 24'b100011001010001110101101;
#10000;
	data_in <= 24'b100101101010110110111000;
#10000;
	data_in <= 24'b110100101101101011011101;
#10000;
	data_in <= 24'b111111111111110011111011;
#10000;
	data_in <= 24'b100011101001110010100011;
#10000;
	data_in <= 24'b010011100110011001110001;
#10000;
	data_in <= 24'b001111000101011001100010;
#10000;
	data_in <= 24'b001110010101001101011111;
#10000;
	data_in <= 24'b001110010101001101011111;
#10000;
	data_in <= 24'b010000000101101001100101;
#10000;
	data_in <= 24'b011001100111101010000010;
#10000;
	data_in <= 24'b110010001100111111010001;
#10000;
	data_in <= 24'b001001010100000101001111;
#10000;
	data_in <= 24'b001011100100100101010110;
#10000;
	data_in <= 24'b001100110100111101011011;
#10000;
	data_in <= 24'b001101000101000001011101;
#10000;
	data_in <= 24'b001101000101000001011101;
#10000;
	data_in <= 24'b001100100100110101011010;
#10000;
	data_in <= 24'b001010000100010001010001;
#10000;
	data_in <= 24'b001100110100111001011010;
#10000;
	data_in <= 24'b001011010100100101010110;
#10000;
	data_in <= 24'b001010110100100001010101;
#10000;
	data_in <= 24'b001010100100011101010100;
#10000;
	data_in <= 24'b001010100100011101010100;
#10000;
	data_in <= 24'b001010100100011101010100;
#10000;
	data_in <= 24'b001010100100011101010101;
#10000;
	data_in <= 24'b001011000100100001010101;
#10000;
	data_in <= 24'b001001100100001001001111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001111101000111010110;
#10000;
	data_in <= 24'b111011001110110011101100;
#10000;
	data_in <= 24'b111110001111011011110101;
#10000;
	data_in <= 24'b111110111111100111111001;
#10000;
	data_in <= 24'b111111001111101111111010;
#10000;
	data_in <= 24'b111110111111101011111001;
#10000;
	data_in <= 24'b111010001110110011101101;
#10000;
	data_in <= 24'b101110001100100111010000;
#10000;
	data_in <= 24'b111101001111000111110001;
#10000;
	data_in <= 24'b111101001111010011110100;
#10000;
	data_in <= 24'b111100101111001011110011;
#10000;
	data_in <= 24'b111100011111001011110010;
#10000;
	data_in <= 24'b111101011111010111110101;
#10000;
	data_in <= 24'b111110011111101011111010;
#10000;
	data_in <= 24'b111111111111111111111110;
#10000;
	data_in <= 24'b111100101111010011110100;
#10000;
	data_in <= 24'b111100111111001011110010;
#10000;
	data_in <= 24'b111011111110111111101111;
#10000;
	data_in <= 24'b111110011111100011111000;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111110011111100111111001;
#10000;
	data_in <= 24'b111110011111101011111010;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111011111111000011110000;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b110001111100100011001011;
#10000;
	data_in <= 24'b011110100111111010000101;
#10000;
	data_in <= 24'b110001111100100111001011;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111110101111101011111010;
#10000;
	data_in <= 24'b111111101111111011111110;
#10000;
	data_in <= 24'b111000101110001111100100;
#10000;
	data_in <= 24'b101100101011010010111000;
#10000;
	data_in <= 24'b100000111000100010001110;
#10000;
	data_in <= 24'b000000100000110100010111;
#10000;
	data_in <= 24'b000111110010011100110000;
#10000;
	data_in <= 24'b101110101011110010111111;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111110111111110011111100;
#10000;
	data_in <= 24'b110011001100110011001100;
#10000;
	data_in <= 24'b001000010010011000101011;
#10000;
	data_in <= 24'b000011010001011100011110;
#10000;
	data_in <= 24'b000011000001100000011111;
#10000;
	data_in <= 24'b000000000000001000001001;
#10000;
	data_in <= 24'b011001100110100001101100;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b111111011111110111111101;
#10000;
	data_in <= 24'b011100101000000110001001;
#10000;
	data_in <= 24'b011111001000011110001101;
#10000;
	data_in <= 24'b011101011000001010001001;
#10000;
	data_in <= 24'b011011000111100010000000;
#10000;
	data_in <= 24'b010001010100111001010101;
#10000;
	data_in <= 24'b100001101000101010001101;
#10000;
	data_in <= 24'b111111101111111011111110;
#10000;
	data_in <= 24'b111111111111111111111111;
#10000;
	data_in <= 24'b000111010011101001001000;
#10000;
	data_in <= 24'b100011001010000010101011;
#10000;
	data_in <= 24'b110110011110011111110000;
#10000;
	data_in <= 24'b110011001101101111100100;
#10000;
	data_in <= 24'b110010101101100111100010;
#10000;
	data_in <= 24'b110001011101001111011100;
#10000;
	data_in <= 24'b110010101101011011011101;
#10000;
	data_in <= 24'b111001001110101011101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000111011101011000100;
#10000;
	data_in <= 24'b101000111011100011000010;
#10000;
	data_in <= 24'b101010101100000011001010;
#10000;
	data_in <= 24'b011001100111110010001001;
#10000;
	data_in <= 24'b000000010001010100100101;
#10000;
	data_in <= 24'b000001010010000000101111;
#10000;
	data_in <= 24'b000001110010000100110000;
#10000;
	data_in <= 24'b000001010001110100101100;
#10000;
	data_in <= 24'b101101001100010111001101;
#10000;
	data_in <= 24'b101000011011011111000010;
#10000;
	data_in <= 24'b101001001011100111000100;
#10000;
	data_in <= 24'b100100111010100110110100;
#10000;
	data_in <= 24'b000110010010111000111101;
#10000;
	data_in <= 24'b000000000001010000100011;
#10000;
	data_in <= 24'b000000100001101100101011;
#10000;
	data_in <= 24'b000000110001101000101001;
#10000;
	data_in <= 24'b110111101110010011100111;
#10000;
	data_in <= 24'b101000111011100111000011;
#10000;
	data_in <= 24'b101000001011010111000000;
#10000;
	data_in <= 24'b101001001011101011000100;
#10000;
	data_in <= 24'b010000010101011001100100;
#10000;
	data_in <= 24'b000000000000111100011111;
#10000;
	data_in <= 24'b000000010001100000101001;
#10000;
	data_in <= 24'b000000100001100000101000;
#10000;
	data_in <= 24'b111101011111011111110111;
#10000;
	data_in <= 24'b101100001100001111001011;
#10000;
	data_in <= 24'b100111111011010010111111;
#10000;
	data_in <= 24'b101001011011101111000100;
#10000;
	data_in <= 24'b011010100111111110001011;
#10000;
	data_in <= 24'b000000000001000100100001;
#10000;
	data_in <= 24'b000000000001010100100110;
#10000;
	data_in <= 24'b000000100001011000100110;
#10000;
	data_in <= 24'b111111001111110011111011;
#10000;
	data_in <= 24'b101110011100100111010001;
#10000;
	data_in <= 24'b100111111011011011000000;
#10000;
	data_in <= 24'b101000111011100011000010;
#10000;
	data_in <= 24'b100001101001110010100111;
#10000;
	data_in <= 24'b000010110001110100101100;
#10000;
	data_in <= 24'b000000000000111100100000;
#10000;
	data_in <= 24'b000000110001010000100100;
#10000;
	data_in <= 24'b111110101111101011111010;
#10000;
	data_in <= 24'b101110001100100111010000;
#10000;
	data_in <= 24'b101000001011011111000001;
#10000;
	data_in <= 24'b101000101011011111000010;
#10000;
	data_in <= 24'b100101011010110010110111;
#10000;
	data_in <= 24'b001000000010110100111100;
#10000;
	data_in <= 24'b000000000000011000010111;
#10000;
	data_in <= 24'b000001000001000100100000;
#10000;
	data_in <= 24'b111110001111100011111000;
#10000;
	data_in <= 24'b101100111100010111001110;
#10000;
	data_in <= 24'b101000101011100111000011;
#10000;
	data_in <= 24'b101000111011100011000010;
#10000;
	data_in <= 24'b100111001011001110111110;
#10000;
	data_in <= 24'b001100110011111001001110;
#10000;
	data_in <= 24'b000000000000000000010000;
#10000;
	data_in <= 24'b000001000000101000011101;
#10000;
	data_in <= 24'b111001101110101011101101;
#10000;
	data_in <= 24'b101010111011111111001001;
#10000;
	data_in <= 24'b101001001011101111000101;
#10000;
	data_in <= 24'b101000111011100011000010;
#10000;
	data_in <= 24'b100111111011011011000001;
#10000;
	data_in <= 24'b010000100100111001011011;
#10000;
	data_in <= 24'b000000010000000100001011;
#10000;
	data_in <= 24'b000000000000000000010011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000000000000111100100000;
#10000;
	data_in <= 24'b010110110101100101001110;
#10000;
	data_in <= 24'b101110111010001001111011;
#10000;
	data_in <= 24'b101100101001101101110110;
#10000;
	data_in <= 24'b101100101001101001110101;
#10000;
	data_in <= 24'b101100011001100001110011;
#10000;
	data_in <= 24'b101100001001011001110001;
#10000;
	data_in <= 24'b101011101001010001101111;
#10000;
	data_in <= 24'b000000000000110000011110;
#10000;
	data_in <= 24'b001111010100000000111110;
#10000;
	data_in <= 24'b101101101001111101111011;
#10000;
	data_in <= 24'b101101101001111101111010;
#10000;
	data_in <= 24'b101101001001110101111000;
#10000;
	data_in <= 24'b101100111001101101110110;
#10000;
	data_in <= 24'b101100101001100101110011;
#10000;
	data_in <= 24'b101100001001011101110001;
#10000;
	data_in <= 24'b000000000000101100011111;
#10000;
	data_in <= 24'b001011010011000100110110;
#10000;
	data_in <= 24'b101011111001101101111001;
#10000;
	data_in <= 24'b101110101010001101111101;
#10000;
	data_in <= 24'b101101101001111101111011;
#10000;
	data_in <= 24'b101101011001110101111001;
#10000;
	data_in <= 24'b101101001001110001110110;
#10000;
	data_in <= 24'b101100101001100101110100;
#10000;
	data_in <= 24'b000000000000101000011101;
#10000;
	data_in <= 24'b001010100010110100110100;
#10000;
	data_in <= 24'b101011101001101001111010;
#10000;
	data_in <= 24'b101111001010010110000000;
#10000;
	data_in <= 24'b101110001010000001111101;
#10000;
	data_in <= 24'b101101111001111101111011;
#10000;
	data_in <= 24'b101101101001111001111000;
#10000;
	data_in <= 24'b101101001001101101110111;
#10000;
	data_in <= 24'b000000000000011000011001;
#10000;
	data_in <= 24'b001100010011001000110101;
#10000;
	data_in <= 24'b101100111001111101111111;
#10000;
	data_in <= 24'b101111011010011010000010;
#10000;
	data_in <= 24'b101110101010001001111111;
#10000;
	data_in <= 24'b101110011010000101111110;
#10000;
	data_in <= 24'b101101111001111101111010;
#10000;
	data_in <= 24'b101101101001110101111001;
#10000;
	data_in <= 24'b000000000000000100010100;
#10000;
	data_in <= 24'b010000100100000000111111;
#10000;
	data_in <= 24'b101111101010100110000101;
#10000;
	data_in <= 24'b101111011010011110000011;
#10000;
	data_in <= 24'b101110111010010110000001;
#10000;
	data_in <= 24'b101110111010001110000000;
#10000;
	data_in <= 24'b101110011010000101111101;
#10000;
	data_in <= 24'b101101111001111101111010;
#10000;
	data_in <= 24'b000000000000000000010010;
#10000;
	data_in <= 24'b011010000101111101010101;
#10000;
	data_in <= 24'b110010011011000110001100;
#10000;
	data_in <= 24'b101111011010011110000100;
#10000;
	data_in <= 24'b101111101010100010000100;
#10000;
	data_in <= 24'b101111001010010110000001;
#10000;
	data_in <= 24'b101110111010001101111110;
#10000;
	data_in <= 24'b101110011010000101111100;
#10000;
	data_in <= 24'b000100110001001000011110;
#10000;
	data_in <= 24'b101001101001010001111010;
#10000;
	data_in <= 24'b110001111011000010001100;
#10000;
	data_in <= 24'b110000001010101010000110;
#10000;
	data_in <= 24'b110000001010100110000110;
#10000;
	data_in <= 24'b101111101010011110000011;
#10000;
	data_in <= 24'b101111001010010110000000;
#10000;
	data_in <= 24'b101110101010001001111110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101011011001001101101101;
#10000;
	data_in <= 24'b101010101001000001101001;
#10000;
	data_in <= 24'b101010001000111001100111;
#10000;
	data_in <= 24'b101001011000101101100101;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b101000011000011101011111;
#10000;
	data_in <= 24'b100111101000010001011100;
#10000;
	data_in <= 24'b100111001000000001011001;
#10000;
	data_in <= 24'b101011101001010101101111;
#10000;
	data_in <= 24'b101011011001010001101101;
#10000;
	data_in <= 24'b101010101001000001101010;
#10000;
	data_in <= 24'b101001111000110101101000;
#10000;
	data_in <= 24'b101001001000101101100101;
#10000;
	data_in <= 24'b101000101000100101100010;
#10000;
	data_in <= 24'b101000001000011101011111;
#10000;
	data_in <= 24'b100111011000001101011100;
#10000;
	data_in <= 24'b101100001001011101110001;
#10000;
	data_in <= 24'b101011101001010101101111;
#10000;
	data_in <= 24'b101011001001001001101101;
#10000;
	data_in <= 24'b101010011000111101101011;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101001001000101101100100;
#10000;
	data_in <= 24'b101000101000100101100001;
#10000;
	data_in <= 24'b100111111000010101011101;
#10000;
	data_in <= 24'b101100101001100101110100;
#10000;
	data_in <= 24'b101100001001011101110001;
#10000;
	data_in <= 24'b101011101001010001101111;
#10000;
	data_in <= 24'b101010111001000101101100;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101001011000110001100110;
#10000;
	data_in <= 24'b101000111000101001100011;
#10000;
	data_in <= 24'b101000001000011001011111;
#10000;
	data_in <= 24'b101101001001101101110110;
#10000;
	data_in <= 24'b101100101001100001110011;
#10000;
	data_in <= 24'b101011111001011001110001;
#10000;
	data_in <= 24'b101011011001001101101110;
#10000;
	data_in <= 24'b101010011001000001101011;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101001011000101101100110;
#10000;
	data_in <= 24'b101000101000100001100010;
#10000;
	data_in <= 24'b101101101001110101111000;
#10000;
	data_in <= 24'b101100111001101101110101;
#10000;
	data_in <= 24'b101100001001100001110010;
#10000;
	data_in <= 24'b101011101001010101110000;
#10000;
	data_in <= 24'b101011001001001101101100;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101000111000100101100100;
#10000;
	data_in <= 24'b101101111001111101111011;
#10000;
	data_in <= 24'b101101011001110101110111;
#10000;
	data_in <= 24'b101100101001101001110100;
#10000;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b101011011001010101101111;
#10000;
	data_in <= 24'b101010101001001001101100;
#10000;
	data_in <= 24'b101001111000111101101000;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101110001010000001111100;
#10000;
	data_in <= 24'b101101111001111001111001;
#10000;
	data_in <= 24'b101101001001101101110110;
#10000;
	data_in <= 24'b101100011001100001110100;
#10000;
	data_in <= 24'b101011101001011001110001;
#10000;
	data_in <= 24'b101010111001001101101101;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100110100111111001010110;
#10000;
	data_in <= 24'b100101110111101101010011;
#10000;
	data_in <= 24'b100101010111100001010000;
#10000;
	data_in <= 24'b100100100111010101001100;
#10000;
	data_in <= 24'b100011110111001001001001;
#10000;
	data_in <= 24'b100010100110111001000101;
#10000;
	data_in <= 24'b100001110110101101000010;
#10000;
	data_in <= 24'b100001000110011100111110;
#10000;
	data_in <= 24'b100110110111111101011000;
#10000;
	data_in <= 24'b100110000111110101010101;
#10000;
	data_in <= 24'b100101100111101001010010;
#10000;
	data_in <= 24'b100100110111011101001110;
#10000;
	data_in <= 24'b100100010111010001001011;
#10000;
	data_in <= 24'b100011000111000001001000;
#10000;
	data_in <= 24'b100010000110110101000100;
#10000;
	data_in <= 24'b100001100110100101000000;
#10000;
	data_in <= 24'b100111001000001001011010;
#10000;
	data_in <= 24'b100110100111111101010111;
#10000;
	data_in <= 24'b100101110111110001010011;
#10000;
	data_in <= 24'b100101000111100101001111;
#10000;
	data_in <= 24'b100100100111010101001101;
#10000;
	data_in <= 24'b100011100111001001001001;
#10000;
	data_in <= 24'b100010010110111001000101;
#10000;
	data_in <= 24'b100001110110101001000010;
#10000;
	data_in <= 24'b100111101000001101011100;
#10000;
	data_in <= 24'b100110111000000001011001;
#10000;
	data_in <= 24'b100110010111111001010110;
#10000;
	data_in <= 24'b100101100111101001010010;
#10000;
	data_in <= 24'b100100110111011001001110;
#10000;
	data_in <= 24'b100011110111001101001011;
#10000;
	data_in <= 24'b100010100110111101000111;
#10000;
	data_in <= 24'b100001110110101101000011;
#10000;
	data_in <= 24'b100111111000010001011111;
#10000;
	data_in <= 24'b100111001000000101011011;
#10000;
	data_in <= 24'b100110100111111101011000;
#10000;
	data_in <= 24'b100101110111110001010100;
#10000;
	data_in <= 24'b100101000111011101010000;
#10000;
	data_in <= 24'b100100000111010001001101;
#10000;
	data_in <= 24'b100010110111000101001001;
#10000;
	data_in <= 24'b100010000110110101000101;
#10000;
	data_in <= 24'b101000011000011101100000;
#10000;
	data_in <= 24'b100111101000010001011100;
#10000;
	data_in <= 24'b100110111000000101011001;
#10000;
	data_in <= 24'b100110000111110101010101;
#10000;
	data_in <= 24'b100101010111101001010001;
#10000;
	data_in <= 24'b100100100111011101001110;
#10000;
	data_in <= 24'b100011010111001101001010;
#10000;
	data_in <= 24'b100010010110111001000110;
#10000;
	data_in <= 24'b101000101000100001100010;
#10000;
	data_in <= 24'b100111111000010101011110;
#10000;
	data_in <= 24'b100111011000001001011011;
#10000;
	data_in <= 24'b100110010111111001010110;
#10000;
	data_in <= 24'b100101100111101101010011;
#10000;
	data_in <= 24'b100100110111100001001111;
#10000;
	data_in <= 24'b100011100111010101001100;
#10000;
	data_in <= 24'b100010100111000001001000;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b101000011000011001100000;
#10000;
	data_in <= 24'b100111101000001101011100;
#10000;
	data_in <= 24'b100110101000000001011000;
#10000;
	data_in <= 24'b100110000111101101010100;
#10000;
	data_in <= 24'b100101000111100101010000;
#10000;
	data_in <= 24'b100011110111010101001101;
#10000;
	data_in <= 24'b100010110111000001001001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100011010111000101001010;
#10000;
	data_in <= 24'b100100010111010101001110;
#10000;
	data_in <= 24'b100101010111101001010010;
#10000;
	data_in <= 24'b100110010111110101010110;
#10000;
	data_in <= 24'b100111001000000101011010;
#10000;
	data_in <= 24'b100111111000010101011110;
#10000;
	data_in <= 24'b101000101000100001100001;
#10000;
	data_in <= 24'b101001011000101001100100;
#10000;
	data_in <= 24'b100011100111001101001011;
#10000;
	data_in <= 24'b100100010111011001001111;
#10000;
	data_in <= 24'b100101100111101101010011;
#10000;
	data_in <= 24'b100110100111111101010111;
#10000;
	data_in <= 24'b100111011000001001011011;
#10000;
	data_in <= 24'b101000001000011001100000;
#10000;
	data_in <= 24'b101000111000100101100010;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
	data_in <= 24'b100011110111010001001101;
#10000;
	data_in <= 24'b100100100111011101010000;
#10000;
	data_in <= 24'b100101100111110001010100;
#10000;
	data_in <= 24'b100110111000000001011001;
#10000;
	data_in <= 24'b100111101000010001011100;
#10000;
	data_in <= 24'b101000011000100001100001;
#10000;
	data_in <= 24'b101001001000101001100100;
#10000;
	data_in <= 24'b101001111000110101101000;
#10000;
	data_in <= 24'b100011110111010001001101;
#10000;
	data_in <= 24'b100100100111100001010001;
#10000;
	data_in <= 24'b100101110111110001010110;
#10000;
	data_in <= 24'b100110111000000001011011;
#10000;
	data_in <= 24'b100111111000010001011101;
#10000;
	data_in <= 24'b101000101000100001100010;
#10000;
	data_in <= 24'b101001011000101101100101;
#10000;
	data_in <= 24'b101010001000111001101010;
#10000;
	data_in <= 24'b100100000111010101001110;
#10000;
	data_in <= 24'b100100110111100101010010;
#10000;
	data_in <= 24'b100101110111111001010111;
#10000;
	data_in <= 24'b100111001000001001011011;
#10000;
	data_in <= 24'b100111111000010101011111;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b101001011000110001100110;
#10000;
	data_in <= 24'b101010011000111101101010;
#10000;
	data_in <= 24'b100100000111011001010000;
#10000;
	data_in <= 24'b100100110111101101010100;
#10000;
	data_in <= 24'b100110001000000001010111;
#10000;
	data_in <= 24'b100111001000001101011100;
#10000;
	data_in <= 24'b101000001000011001100000;
#10000;
	data_in <= 24'b101001001000101001100100;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101010011001000001101100;
#10000;
	data_in <= 24'b100100010111011001010000;
#10000;
	data_in <= 24'b100101000111101101010100;
#10000;
	data_in <= 24'b100110001000000001011000;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b101000011000011101100001;
#10000;
	data_in <= 24'b101001001000101001100101;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b100100010111011101010001;
#10000;
	data_in <= 24'b100101000111101101010101;
#10000;
	data_in <= 24'b100110011000000101011001;
#10000;
	data_in <= 24'b100111101000010001011110;
#10000;
	data_in <= 24'b101000101000011101100010;
#10000;
	data_in <= 24'b101001011000101101100110;
#10000;
	data_in <= 24'b101010001000111101101001;
#10000;
	data_in <= 24'b101010111001001001101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101010001000111001101000;
#10000;
	data_in <= 24'b101010111001001001101100;
#10000;
	data_in <= 24'b101011011001010101101111;
#10000;
	data_in <= 24'b101100001001011101110010;
#10000;
	data_in <= 24'b101101001001101001110110;
#10000;
	data_in <= 24'b101101111001110001111000;
#10000;
	data_in <= 24'b101110011010000001111010;
#10000;
	data_in <= 24'b101110111010001001111110;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101011001001010001101101;
#10000;
	data_in <= 24'b101011101001011001110000;
#10000;
	data_in <= 24'b101100011001100001110100;
#10000;
	data_in <= 24'b101101011001101101110111;
#10000;
	data_in <= 24'b101101111001111101111010;
#10000;
	data_in <= 24'b101110101010001001111100;
#10000;
	data_in <= 24'b101111001010010001111111;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101011011001010101101111;
#10000;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b101100101001101001110101;
#10000;
	data_in <= 24'b101101101001110101111001;
#10000;
	data_in <= 24'b101110011001111101111011;
#10000;
	data_in <= 24'b101110111010001001111110;
#10000;
	data_in <= 24'b101111011010010110000001;
#10000;
	data_in <= 24'b101010111001001001101101;
#10000;
	data_in <= 24'b101011011001011001110000;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b101100111001101101110110;
#10000;
	data_in <= 24'b101101111001110101111001;
#10000;
	data_in <= 24'b101110101010000001111101;
#10000;
	data_in <= 24'b101111001010001110000000;
#10000;
	data_in <= 24'b101111101010011010000011;
#10000;
	data_in <= 24'b101011001001001101101110;
#10000;
	data_in <= 24'b101011101001011101110001;
#10000;
	data_in <= 24'b101100011001101001110100;
#10000;
	data_in <= 24'b101101001001110001110111;
#10000;
	data_in <= 24'b101110001001111101111011;
#10000;
	data_in <= 24'b101110111010001101111101;
#10000;
	data_in <= 24'b101111001010010110000000;
#10000;
	data_in <= 24'b101111111010100010000100;
#10000;
	data_in <= 24'b101011011001010001110000;
#10000;
	data_in <= 24'b101011111001100001110010;
#10000;
	data_in <= 24'b101100101001101101110101;
#10000;
	data_in <= 24'b101101011001111001111001;
#10000;
	data_in <= 24'b101110001010000101111100;
#10000;
	data_in <= 24'b101110111010010001111111;
#10000;
	data_in <= 24'b101111101010011110000010;
#10000;
	data_in <= 24'b110000001010100110000101;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b101100101001101101110110;
#10000;
	data_in <= 24'b101101101001111001111010;
#10000;
	data_in <= 24'b101110011010000101111101;
#10000;
	data_in <= 24'b101111001010010110000000;
#10000;
	data_in <= 24'b101111101010011110000011;
#10000;
	data_in <= 24'b110000011010101010000110;
#10000;
	data_in <= 24'b101011101001010101110001;
#10000;
	data_in <= 24'b101100001001100101110100;
#10000;
	data_in <= 24'b101100111001110001111000;
#10000;
	data_in <= 24'b101101111001111101111100;
#10000;
	data_in <= 24'b101110101010001001111110;
#10000;
	data_in <= 24'b101111011010011010000001;
#10000;
	data_in <= 24'b101111111010100010000101;
#10000;
	data_in <= 24'b110000011010101010000111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101111001010001110000000;
#10000;
	data_in <= 24'b101111101010011010000010;
#10000;
	data_in <= 24'b110000011010100110000101;
#10000;
	data_in <= 24'b110000101010101110001000;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110001011010111010001011;
#10000;
	data_in <= 24'b110001101010111110001100;
#10000;
	data_in <= 24'b110010011011001010001111;
#10000;
	data_in <= 24'b101111101010011010000010;
#10000;
	data_in <= 24'b110000001010100010000100;
#10000;
	data_in <= 24'b110000011010101010000111;
#10000;
	data_in <= 24'b110000111010110110001010;
#10000;
	data_in <= 24'b110001011010111110001011;
#10000;
	data_in <= 24'b110001101011000010001100;
#10000;
	data_in <= 24'b110010011011001010001111;
#10000;
	data_in <= 24'b110010111011010010010001;
#10000;
	data_in <= 24'b101111111010011110000100;
#10000;
	data_in <= 24'b110000011010100110000101;
#10000;
	data_in <= 24'b110000101010101110001000;
#10000;
	data_in <= 24'b110001011010111010001011;
#10000;
	data_in <= 24'b110001101011000010001100;
#10000;
	data_in <= 24'b110001111011000110001110;
#10000;
	data_in <= 24'b110010101011001110010001;
#10000;
	data_in <= 24'b110011001011010110010011;
#10000;
	data_in <= 24'b110000001010100010000101;
#10000;
	data_in <= 24'b110000101010101010000111;
#10000;
	data_in <= 24'b110001001010110110001001;
#10000;
	data_in <= 24'b110001011010111010001011;
#10000;
	data_in <= 24'b110001111011000110001110;
#10000;
	data_in <= 24'b110010011011001110010000;
#10000;
	data_in <= 24'b110010111011010010010010;
#10000;
	data_in <= 24'b110011101011011010010100;
#10000;
	data_in <= 24'b110000011010100110000110;
#10000;
	data_in <= 24'b110000111010101110001000;
#10000;
	data_in <= 24'b110001011010111010001010;
#10000;
	data_in <= 24'b110001101011000110001101;
#10000;
	data_in <= 24'b110010001011001110010000;
#10000;
	data_in <= 24'b110010011011010010010001;
#10000;
	data_in <= 24'b110011001011011010010011;
#10000;
	data_in <= 24'b110011111011011110010110;
#10000;
	data_in <= 24'b110000101010101110000111;
#10000;
	data_in <= 24'b110001001010110110001010;
#10000;
	data_in <= 24'b110001011010111110001100;
#10000;
	data_in <= 24'b110001111011001010001111;
#10000;
	data_in <= 24'b110010011011010010010010;
#10000;
	data_in <= 24'b110010101011010110010011;
#10000;
	data_in <= 24'b110011011011011110010110;
#10000;
	data_in <= 24'b110011111011100010010111;
#10000;
	data_in <= 24'b110000111010101110001000;
#10000;
	data_in <= 24'b110001011010111010001010;
#10000;
	data_in <= 24'b110001101011000010001101;
#10000;
	data_in <= 24'b110010001011001110010000;
#10000;
	data_in <= 24'b110010101011010110010010;
#10000;
	data_in <= 24'b110010111011011110010101;
#10000;
	data_in <= 24'b110011101011100010010110;
#10000;
	data_in <= 24'b110100001011100110011000;
#10000;
	data_in <= 24'b110000111010110010001010;
#10000;
	data_in <= 24'b110001011010111010001100;
#10000;
	data_in <= 24'b110001111011000110001111;
#10000;
	data_in <= 24'b110010011011010010010010;
#10000;
	data_in <= 24'b110010101011011010010100;
#10000;
	data_in <= 24'b110011001011011110010110;
#10000;
	data_in <= 24'b110011111011100010010111;
#10000;
	data_in <= 24'b110100011011101010011001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110010111011001110010001;
#10000;
	data_in <= 24'b110011001011010010010010;
#10000;
	data_in <= 24'b110011011011011010010011;
#10000;
	data_in <= 24'b110011011011011010010101;
#10000;
	data_in <= 24'b110011011011011110010110;
#10000;
	data_in <= 24'b110011111011100110011000;
#10000;
	data_in <= 24'b110001011011000110010011;
#10000;
	data_in <= 24'b010010010100010001000011;
#10000;
	data_in <= 24'b110011001011010110010010;
#10000;
	data_in <= 24'b110011011011011110010011;
#10000;
	data_in <= 24'b110011101011100010010101;
#10000;
	data_in <= 24'b110011111011100110010111;
#10000;
	data_in <= 24'b110011111011101010011000;
#10000;
	data_in <= 24'b110011111011100110011000;
#10000;
	data_in <= 24'b110100011011110010011011;
#10000;
	data_in <= 24'b110001101011010010010110;
#10000;
	data_in <= 24'b110011011011011110010100;
#10000;
	data_in <= 24'b110011101011100010010101;
#10000;
	data_in <= 24'b110011111011100110010111;
#10000;
	data_in <= 24'b110100001011101010011001;
#10000;
	data_in <= 24'b110100011011101110011010;
#10000;
	data_in <= 24'b110100101011110010011011;
#10000;
	data_in <= 24'b110100001011101110011011;
#10000;
	data_in <= 24'b110101001011111110011110;
#10000;
	data_in <= 24'b110011111011100010010110;
#10000;
	data_in <= 24'b110011111011100110010111;
#10000;
	data_in <= 24'b110100001011101010011001;
#10000;
	data_in <= 24'b110100011011101110011010;
#10000;
	data_in <= 24'b110100101011110010011100;
#10000;
	data_in <= 24'b110100111011110110011101;
#10000;
	data_in <= 24'b110101001011111010011101;
#10000;
	data_in <= 24'b110101001011111110011110;
#10000;
	data_in <= 24'b110011111011100110010111;
#10000;
	data_in <= 24'b110100001011101110011000;
#10000;
	data_in <= 24'b110100101011110010011011;
#10000;
	data_in <= 24'b110100111011110110011100;
#10000;
	data_in <= 24'b110100111011111010011101;
#10000;
	data_in <= 24'b110101001011111110011111;
#10000;
	data_in <= 24'b110101011100000010011111;
#10000;
	data_in <= 24'b110101011100000010011111;
#10000;
	data_in <= 24'b110100001011101010011000;
#10000;
	data_in <= 24'b110100101011110110011011;
#10000;
	data_in <= 24'b110100111011111010011100;
#10000;
	data_in <= 24'b110101001011111110011101;
#10000;
	data_in <= 24'b110101001100000010011111;
#10000;
	data_in <= 24'b110101011100000010100000;
#10000;
	data_in <= 24'b110101011100000010100000;
#10000;
	data_in <= 24'b110101111100001010100010;
#10000;
	data_in <= 24'b110100011011101110011010;
#10000;
	data_in <= 24'b110100111011111010011100;
#10000;
	data_in <= 24'b110100111011111010011101;
#10000;
	data_in <= 24'b110101011100000010011110;
#10000;
	data_in <= 24'b110101011100000010100000;
#10000;
	data_in <= 24'b110101101100000110100001;
#10000;
	data_in <= 24'b110101101100000110100001;
#10000;
	data_in <= 24'b110101111100001110100010;
#10000;
	data_in <= 24'b110100101011110010011011;
#10000;
	data_in <= 24'b110101001011111110011110;
#10000;
	data_in <= 24'b110101011100000010011110;
#10000;
	data_in <= 24'b110101011100000010011111;
#10000;
	data_in <= 24'b110101101100000110100001;
#10000;
	data_in <= 24'b110101111100001010100010;
#10000;
	data_in <= 24'b110101111100001010100011;
#10000;
	data_in <= 24'b110110011100010010100100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000000000000000000000000;
#10000;
	data_in <= 24'b000101010001101000101011;
#10000;
	data_in <= 24'b100100111010101010110101;
#10000;
	data_in <= 24'b101000111011100111000011;
#10000;
	data_in <= 24'b101001101011101111000100;
#10000;
	data_in <= 24'b101001101011110011000110;
#10000;
	data_in <= 24'b101100011100001111001011;
#10000;
	data_in <= 24'b110010111101010111011011;
#10000;
	data_in <= 24'b011010110110000101010110;
#10000;
	data_in <= 24'b010000100100010101001100;
#10000;
	data_in <= 24'b100100111010101010110101;
#10000;
	data_in <= 24'b101000111011100011000010;
#10000;
	data_in <= 24'b101001001011101011000011;
#10000;
	data_in <= 24'b101100011100001111001100;
#10000;
	data_in <= 24'b101111111100111011010111;
#10000;
	data_in <= 24'b110000111101001111011100;
#10000;
	data_in <= 24'b110101101100000110011110;
#10000;
	data_in <= 24'b101011101010100110010111;
#10000;
	data_in <= 24'b100011111010100010110011;
#10000;
	data_in <= 24'b101000001011011011000000;
#10000;
	data_in <= 24'b101100101100001111001101;
#10000;
	data_in <= 24'b110001001101001011011011;
#10000;
	data_in <= 24'b110010011101100011100000;
#10000;
	data_in <= 24'b110011001101101111100011;
#10000;
	data_in <= 24'b110101001011111010011100;
#10000;
	data_in <= 24'b101101011010110110011001;
#10000;
	data_in <= 24'b100010111010001110101110;
#10000;
	data_in <= 24'b101011101100000011001001;
#10000;
	data_in <= 24'b110001101101010011011100;
#10000;
	data_in <= 24'b110010011101100011100000;
#10000;
	data_in <= 24'b110011011101110011100100;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110110001100001010011111;
#10000;
	data_in <= 24'b101110001010110110010111;
#10000;
	data_in <= 24'b100110011010110010110100;
#10000;
	data_in <= 24'b110001001101001111011011;
#10000;
	data_in <= 24'b110010101101100111100000;
#10000;
	data_in <= 24'b110011101101110111100100;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110101111100001010100000;
#10000;
	data_in <= 24'b110000101011010110011101;
#10000;
	data_in <= 24'b101110001100011011001100;
#10000;
	data_in <= 24'b110010011101100111100010;
#10000;
	data_in <= 24'b110011011101101111100011;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110110001100000110100000;
#10000;
	data_in <= 24'b110001101100000110110010;
#10000;
	data_in <= 24'b110001001101010011011110;
#10000;
	data_in <= 24'b110011001101101011100010;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110101101100000110100001;
#10000;
	data_in <= 24'b110000101100101011001000;
#10000;
	data_in <= 24'b110001111101011111100001;
#10000;
	data_in <= 24'b110011101101110011100011;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110000101101000111011001;
#10000;
	data_in <= 24'b110000011101000111011010;
#10000;
	data_in <= 24'b110011001101110011100100;
#10000;
	data_in <= 24'b110011001101101111100011;
#10000;
	data_in <= 24'b110101001110001111101011;
#10000;
	data_in <= 24'b011111001001000010011011;
#10000;
	data_in <= 24'b000011010010101000111001;
#10000;
	data_in <= 24'b000111110011110001001010;
#10000;
	data_in <= 24'b110010011101100011100000;
#10000;
	data_in <= 24'b110011001101101111100011;
#10000;
	data_in <= 24'b110011001101101111100011;
#10000;
	data_in <= 24'b110011011101110011100100;
#10000;
	data_in <= 24'b110101101110010011101100;
#10000;
	data_in <= 24'b010101110110111001111010;
#10000;
	data_in <= 24'b000000010001111100101110;
#10000;
	data_in <= 24'b000100010010111100111110;
#10000;
	data_in <= 24'b110011101101110011100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110101101110010111101101;
#10000;
	data_in <= 24'b010100110110100001110100;
#10000;
	data_in <= 24'b000000010001010100100101;
#10000;
	data_in <= 24'b000001100010010100110101;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110110011110100011101111;
#10000;
	data_in <= 24'b011101001000011110010011;
#10000;
	data_in <= 24'b000000000000111000011101;
#10000;
	data_in <= 24'b000000100010000100110000;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110101001110001111101010;
#10000;
	data_in <= 24'b101110111100110111010100;
#10000;
	data_in <= 24'b001100000100011101010101;
#10000;
	data_in <= 24'b000000000001001000100001;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110101001110001011101010;
#10000;
	data_in <= 24'b101110111100110011010100;
#10000;
	data_in <= 24'b011110001000101110010110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110100111110001011101001;
#10000;
	data_in <= 24'b110110001110011111101110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000111000011101001001000;
#10000;
	data_in <= 24'b000111000011101001001001;
#10000;
	data_in <= 24'b000111000011101001001001;
#10000;
	data_in <= 24'b000111000011101001001001;
#10000;
	data_in <= 24'b000111000011101001001001;
#10000;
	data_in <= 24'b000111000011101001001001;
#10000;
	data_in <= 24'b000111000011101001001001;
#10000;
	data_in <= 24'b000111110011110001001010;
#10000;
	data_in <= 24'b000011100010110100111100;
#10000;
	data_in <= 24'b000011110010110100111100;
#10000;
	data_in <= 24'b000011110010110100111100;
#10000;
	data_in <= 24'b000011110010110100111100;
#10000;
	data_in <= 24'b000011110010110100111100;
#10000;
	data_in <= 24'b000011110010110100111100;
#10000;
	data_in <= 24'b000011110010110100111101;
#10000;
	data_in <= 24'b000100000010111000111101;
#10000;
	data_in <= 24'b000001000010001100110011;
#10000;
	data_in <= 24'b000001000010001100110011;
#10000;
	data_in <= 24'b000001000010001100110011;
#10000;
	data_in <= 24'b000001000010010000110011;
#10000;
	data_in <= 24'b000001000010010000110011;
#10000;
	data_in <= 24'b000001000010001100110011;
#10000;
	data_in <= 24'b000001000010001100110011;
#10000;
	data_in <= 24'b000001010010010000110100;
#10000;
	data_in <= 24'b000000010010000100110000;
#10000;
	data_in <= 24'b000000000010000000110000;
#10000;
	data_in <= 24'b000000000001111100101111;
#10000;
	data_in <= 24'b000000000001110000101011;
#10000;
	data_in <= 24'b000000000001110000101011;
#10000;
	data_in <= 24'b000000000001111100101110;
#10000;
	data_in <= 24'b000000000001111100101110;
#10000;
	data_in <= 24'b000000000001111100101111;
#10000;
	data_in <= 24'b000000000001011000100110;
#10000;
	data_in <= 24'b000000000001010100100101;
#10000;
	data_in <= 24'b000000000001101000101001;
#10000;
	data_in <= 24'b000100100010110100111101;
#10000;
	data_in <= 24'b000100000010110000111011;
#10000;
	data_in <= 24'b000000000001110100101100;
#10000;
	data_in <= 24'b000000000001101000101001;
#10000;
	data_in <= 24'b000000010001110100101100;
#10000;
	data_in <= 24'b010110100111000001111011;
#10000;
	data_in <= 24'b011000110111100010000011;
#10000;
	data_in <= 24'b100001011001100010100010;
#10000;
	data_in <= 24'b101011111100000011001001;
#10000;
	data_in <= 24'b101011011011111011000110;
#10000;
	data_in <= 24'b100100101010010110101110;
#10000;
	data_in <= 24'b100010011001101110100110;
#10000;
	data_in <= 24'b100101101010100110110010;
#10000;
	data_in <= 24'b110101101110010111101100;
#10000;
	data_in <= 24'b110101111110011011101101;
#10000;
	data_in <= 24'b110110001110011111101110;
#10000;
	data_in <= 24'b110101011110010011101011;
#10000;
	data_in <= 24'b110101011110010011101011;
#10000;
	data_in <= 24'b110110001110011111101101;
#10000;
	data_in <= 24'b110110011110011111101110;
#10000;
	data_in <= 24'b110110001110011011101101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000101000011000100111111;
#10000;
	data_in <= 24'b001100000100101101010111;
#10000;
	data_in <= 24'b110000011101000011011000;
#10000;
	data_in <= 24'b110011101101110011100100;
#10000;
	data_in <= 24'b110010011101100011100000;
#10000;
	data_in <= 24'b110010101101100111100001;
#10000;
	data_in <= 24'b110000111101001111011100;
#10000;
	data_in <= 24'b110000011101000011011001;
#10000;
	data_in <= 24'b000010110010100100110111;
#10000;
	data_in <= 24'b000100110011000000111110;
#10000;
	data_in <= 24'b101001111011100011000001;
#10000;
	data_in <= 24'b110110011110011111101111;
#10000;
	data_in <= 24'b110010111101101111100011;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011011101110011100100;
#10000;
	data_in <= 24'b110010111101101011100010;
#10000;
	data_in <= 24'b000000100010000000101111;
#10000;
	data_in <= 24'b000011010010011100110101;
#10000;
	data_in <= 24'b101001111011100111000010;
#10000;
	data_in <= 24'b110110011110011111101111;
#10000;
	data_in <= 24'b110011001101101111100100;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b000000000000111100011111;
#10000;
	data_in <= 24'b001010100100001001001111;
#10000;
	data_in <= 24'b110001111101011111011111;
#10000;
	data_in <= 24'b110100101110000011101000;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b001010010011111001001100;
#10000;
	data_in <= 24'b100111101011000010111001;
#10000;
	data_in <= 24'b110101101110010111101100;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b101111101100111111010111;
#10000;
	data_in <= 24'b110101001110001111101011;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100111110001011101001;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110000011100111111010111;
#10000;
	data_in <= 24'b101011111100001011001011;
#10000;
	data_in <= 24'b101001011011101111000100;
#10000;
	data_in <= 24'b101000111011100011000010;
#10000;
	data_in <= 24'b101000011011100111000011;
#10000;
	data_in <= 24'b010010100101100001100011;
#10000;
	data_in <= 24'b000000000000000000000000;
#10000;
	data_in <= 24'b000001110000011100010011;
#10000;
	data_in <= 24'b110001101101011011011110;
#10000;
	data_in <= 24'b110000101101000111011010;
#10000;
	data_in <= 24'b101100101100010011001101;
#10000;
	data_in <= 24'b101000011011011011000000;
#10000;
	data_in <= 24'b100111111011011111000001;
#10000;
	data_in <= 24'b010111010110101001110010;
#10000;
	data_in <= 24'b001110100011010000101110;
#10000;
	data_in <= 24'b100100001000001101101111;
#10000;
	data_in <= 24'b110011001101101111100100;
#10000;
	data_in <= 24'b110010001101011111100000;
#10000;
	data_in <= 24'b110001011101010011011100;
#10000;
	data_in <= 24'b101100101100001111001100;
#10000;
	data_in <= 24'b100101001010110110111001;
#10000;
	data_in <= 24'b100101101001111110011011;
#10000;
	data_in <= 24'b110001001010111110001101;
#10000;
	data_in <= 24'b110100011011101110011000;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011011101110011100100;
#10000;
	data_in <= 24'b110010011101100111100000;
#10000;
	data_in <= 24'b110001111101010111011100;
#10000;
	data_in <= 24'b101000011011011111000011;
#10000;
	data_in <= 24'b100110011010000010011001;
#10000;
	data_in <= 24'b110010111011010110010010;
#10000;
	data_in <= 24'b110011011011011110010110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011101101110111100100;
#10000;
	data_in <= 24'b110010111101100111100000;
#10000;
	data_in <= 24'b101111011100111011011000;
#10000;
	data_in <= 24'b101010101010101010100000;
#10000;
	data_in <= 24'b110011001011011010010010;
#10000;
	data_in <= 24'b110100001011101010011000;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011011101101111100010;
#10000;
	data_in <= 24'b110001111101011111100001;
#10000;
	data_in <= 24'b101111111100001110111110;
#10000;
	data_in <= 24'b110010101011011010010011;
#10000;
	data_in <= 24'b110100011011101110011010;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110011101101110111100100;
#10000;
	data_in <= 24'b110010101101101011100010;
#10000;
	data_in <= 24'b110000011100111111010101;
#10000;
	data_in <= 24'b110010011011101110100010;
#10000;
	data_in <= 24'b110100101011101110010111;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110011111101111111100101;
#10000;
	data_in <= 24'b110011011101110011100001;
#10000;
	data_in <= 24'b110000111101010011011110;
#10000;
	data_in <= 24'b110001011100000110110011;
#10000;
	data_in <= 24'b110100111011101010010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011110010110110101100000;
#10000;
	data_in <= 24'b110010101011001110010000;
#10000;
	data_in <= 24'b110000101010101110001001;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110000101010101110001000;
#10000;
	data_in <= 24'b110000011010100110000101;
#10000;
	data_in <= 24'b101111101010011010000010;
#10000;
	data_in <= 24'b101111001010001110000000;
#10000;
	data_in <= 24'b110010111011010010010010;
#10000;
	data_in <= 24'b110001111011000010001110;
#10000;
	data_in <= 24'b110001101011000010001100;
#10000;
	data_in <= 24'b110001011010111110001011;
#10000;
	data_in <= 24'b110000111010110110001010;
#10000;
	data_in <= 24'b110000011010101010000111;
#10000;
	data_in <= 24'b110000001010100010000100;
#10000;
	data_in <= 24'b101111101010011010000010;
#10000;
	data_in <= 24'b110010111011010010010010;
#10000;
	data_in <= 24'b110010101011001110010000;
#10000;
	data_in <= 24'b110001111011000110001110;
#10000;
	data_in <= 24'b110001101011000010001100;
#10000;
	data_in <= 24'b110001011010111010001011;
#10000;
	data_in <= 24'b110000101010101110001000;
#10000;
	data_in <= 24'b110000011010100110000101;
#10000;
	data_in <= 24'b101111111010011110000100;
#10000;
	data_in <= 24'b110011011011011010010100;
#10000;
	data_in <= 24'b110010111011010010010010;
#10000;
	data_in <= 24'b110010011011001110010000;
#10000;
	data_in <= 24'b110001111011000110001110;
#10000;
	data_in <= 24'b110001011010111010001011;
#10000;
	data_in <= 24'b110001001010110110001001;
#10000;
	data_in <= 24'b110000101010101010000111;
#10000;
	data_in <= 24'b110000001010100010000101;
#10000;
	data_in <= 24'b110011111011100010010110;
#10000;
	data_in <= 24'b110011001011011010010011;
#10000;
	data_in <= 24'b110010011011010010010001;
#10000;
	data_in <= 24'b110010001011001110010000;
#10000;
	data_in <= 24'b110001101011000110001101;
#10000;
	data_in <= 24'b110001011010111010001010;
#10000;
	data_in <= 24'b110000111010101110001000;
#10000;
	data_in <= 24'b110000011010100110000110;
#10000;
	data_in <= 24'b110011111011100010010111;
#10000;
	data_in <= 24'b110011011011011110010110;
#10000;
	data_in <= 24'b110010101011010110010011;
#10000;
	data_in <= 24'b110010011011010010010010;
#10000;
	data_in <= 24'b110001111011001010001111;
#10000;
	data_in <= 24'b110001011010111110001100;
#10000;
	data_in <= 24'b110001001010110110001010;
#10000;
	data_in <= 24'b110000101010101110000111;
#10000;
	data_in <= 24'b110100001011100110011001;
#10000;
	data_in <= 24'b110011101011100010010110;
#10000;
	data_in <= 24'b110010111011011110010101;
#10000;
	data_in <= 24'b110010101011010110010010;
#10000;
	data_in <= 24'b110010001011001110010000;
#10000;
	data_in <= 24'b110001101011000010001101;
#10000;
	data_in <= 24'b110001011010111010001010;
#10000;
	data_in <= 24'b110000111010101110001000;
#10000;
	data_in <= 24'b110100011011101010011010;
#10000;
	data_in <= 24'b110011111011100010010111;
#10000;
	data_in <= 24'b110011001011011110010110;
#10000;
	data_in <= 24'b110010101011011010010100;
#10000;
	data_in <= 24'b110010011011010010010010;
#10000;
	data_in <= 24'b110001111011000110001111;
#10000;
	data_in <= 24'b110001011010111010001100;
#10000;
	data_in <= 24'b110000111010110010001010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101110111010001001111110;
#10000;
	data_in <= 24'b101110011010000001111010;
#10000;
	data_in <= 24'b101101111001110001111000;
#10000;
	data_in <= 24'b101101001001101001110110;
#10000;
	data_in <= 24'b101100001001011101110010;
#10000;
	data_in <= 24'b101011011001010101101111;
#10000;
	data_in <= 24'b101010111001001001101100;
#10000;
	data_in <= 24'b101010001000111001101000;
#10000;
	data_in <= 24'b101111001010010001111111;
#10000;
	data_in <= 24'b101110101010001001111100;
#10000;
	data_in <= 24'b101101111001111101111010;
#10000;
	data_in <= 24'b101101011001101101110111;
#10000;
	data_in <= 24'b101100011001100001110100;
#10000;
	data_in <= 24'b101011101001011001110000;
#10000;
	data_in <= 24'b101011001001010001101101;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101111011010010110000001;
#10000;
	data_in <= 24'b101110111010001001111110;
#10000;
	data_in <= 24'b101110011001111101111011;
#10000;
	data_in <= 24'b101101101001110101111001;
#10000;
	data_in <= 24'b101100101001101001110101;
#10000;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b101011011001010101101111;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101111101010011010000011;
#10000;
	data_in <= 24'b101111001010001110000000;
#10000;
	data_in <= 24'b101110101010000001111101;
#10000;
	data_in <= 24'b101101111001110101111001;
#10000;
	data_in <= 24'b101100111001101101110110;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b101011011001011001110000;
#10000;
	data_in <= 24'b101010111001001001101101;
#10000;
	data_in <= 24'b101111111010100010000100;
#10000;
	data_in <= 24'b101111001010010110000000;
#10000;
	data_in <= 24'b101110111010001101111101;
#10000;
	data_in <= 24'b101110001001111101111011;
#10000;
	data_in <= 24'b101101001001110001110111;
#10000;
	data_in <= 24'b101100011001101001110100;
#10000;
	data_in <= 24'b101011101001011101110001;
#10000;
	data_in <= 24'b101011001001001101101110;
#10000;
	data_in <= 24'b110000001010100110000101;
#10000;
	data_in <= 24'b101111101010011110000010;
#10000;
	data_in <= 24'b101110111010010001111111;
#10000;
	data_in <= 24'b101110001010000101111100;
#10000;
	data_in <= 24'b101101011001111001111001;
#10000;
	data_in <= 24'b101100101001101101110101;
#10000;
	data_in <= 24'b101011111001100001110010;
#10000;
	data_in <= 24'b101011011001010001110000;
#10000;
	data_in <= 24'b110000011010101010000110;
#10000;
	data_in <= 24'b101111101010011110000011;
#10000;
	data_in <= 24'b101111001010010110000000;
#10000;
	data_in <= 24'b101110011010000101111101;
#10000;
	data_in <= 24'b101101101001111001111010;
#10000;
	data_in <= 24'b101100101001101101110110;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b110000011010101010000111;
#10000;
	data_in <= 24'b101111111010100010000101;
#10000;
	data_in <= 24'b101111011010011010000001;
#10000;
	data_in <= 24'b101110101010001001111110;
#10000;
	data_in <= 24'b101101111001111101111100;
#10000;
	data_in <= 24'b101100111001110001111000;
#10000;
	data_in <= 24'b101100001001100101110100;
#10000;
	data_in <= 24'b101011101001010101110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101001011000101001100100;
#10000;
	data_in <= 24'b101000101000100001100001;
#10000;
	data_in <= 24'b100111111000010101011110;
#10000;
	data_in <= 24'b100111001000000101011010;
#10000;
	data_in <= 24'b100110010111110101010110;
#10000;
	data_in <= 24'b100101010111101001010010;
#10000;
	data_in <= 24'b100100010111010101001110;
#10000;
	data_in <= 24'b100011010111000101001010;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
	data_in <= 24'b101000111000100101100010;
#10000;
	data_in <= 24'b101000001000011001100000;
#10000;
	data_in <= 24'b100111011000001001011011;
#10000;
	data_in <= 24'b100110100111111101010111;
#10000;
	data_in <= 24'b100101100111101101010011;
#10000;
	data_in <= 24'b100100010111011001001111;
#10000;
	data_in <= 24'b100011100111001101001011;
#10000;
	data_in <= 24'b101001111000110101101000;
#10000;
	data_in <= 24'b101001001000101001100100;
#10000;
	data_in <= 24'b101000011000100001100001;
#10000;
	data_in <= 24'b100111101000010001011100;
#10000;
	data_in <= 24'b100110111000000001011001;
#10000;
	data_in <= 24'b100101100111110001010100;
#10000;
	data_in <= 24'b100100100111011101010000;
#10000;
	data_in <= 24'b100011110111010001001101;
#10000;
	data_in <= 24'b101010001000111001101010;
#10000;
	data_in <= 24'b101001011000101101100101;
#10000;
	data_in <= 24'b101000101000100001100010;
#10000;
	data_in <= 24'b100111111000010001011101;
#10000;
	data_in <= 24'b100110111000000001011011;
#10000;
	data_in <= 24'b100101110111110001010110;
#10000;
	data_in <= 24'b100100100111100001010001;
#10000;
	data_in <= 24'b100011110111010001001101;
#10000;
	data_in <= 24'b101010011000111101101010;
#10000;
	data_in <= 24'b101001011000110001100110;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b100111111000010101011111;
#10000;
	data_in <= 24'b100111001000001001011011;
#10000;
	data_in <= 24'b100101110111111001010111;
#10000;
	data_in <= 24'b100100110111100101010010;
#10000;
	data_in <= 24'b100100000111010101001110;
#10000;
	data_in <= 24'b101010011001000001101100;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101001001000101001100100;
#10000;
	data_in <= 24'b101000001000011001100000;
#10000;
	data_in <= 24'b100111001000001101011100;
#10000;
	data_in <= 24'b100110001000000001010111;
#10000;
	data_in <= 24'b100100110111101101010100;
#10000;
	data_in <= 24'b100100000111011001010000;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101001001000101001100101;
#10000;
	data_in <= 24'b101000011000011101100001;
#10000;
	data_in <= 24'b100111011000001101011101;
#10000;
	data_in <= 24'b100110001000000001011000;
#10000;
	data_in <= 24'b100101000111101101010100;
#10000;
	data_in <= 24'b100100010111011001010000;
#10000;
	data_in <= 24'b101010111001001001101101;
#10000;
	data_in <= 24'b101010001000111101101001;
#10000;
	data_in <= 24'b101001011000101101100110;
#10000;
	data_in <= 24'b101000101000011101100010;
#10000;
	data_in <= 24'b100111101000010001011110;
#10000;
	data_in <= 24'b100110011000000101011001;
#10000;
	data_in <= 24'b100101000111101101010101;
#10000;
	data_in <= 24'b100100010111011101010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b100101100111110101010110;
#10000;
	data_in <= 24'b100110101000001001011001;
#10000;
	data_in <= 24'b100111101000010101011110;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101011001001001101101110;
#10000;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b100101110111111001010111;
#10000;
	data_in <= 24'b100110101000001001011011;
#10000;
	data_in <= 24'b100111111000011001011111;
#10000;
	data_in <= 24'b101000111000100101100100;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101010011001000001101011;
#10000;
	data_in <= 24'b101011011001010001101111;
#10000;
	data_in <= 24'b100100110111100101010010;
#10000;
	data_in <= 24'b100101100111111001010111;
#10000;
	data_in <= 24'b100110111000001101011100;
#10000;
	data_in <= 24'b100111111000010101100000;
#10000;
	data_in <= 24'b101001001000100101100101;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101010101001000001101011;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b100100110111101001010011;
#10000;
	data_in <= 24'b100101110111111001011000;
#10000;
	data_in <= 24'b100110111000001101011101;
#10000;
	data_in <= 24'b100111111000011001100001;
#10000;
	data_in <= 24'b101001001000101001100101;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b100100110111101101010100;
#10000;
	data_in <= 24'b100101110111111101011000;
#10000;
	data_in <= 24'b100110111000010001011110;
#10000;
	data_in <= 24'b100111111000011101100001;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101010101001001001101101;
#10000;
	data_in <= 24'b101011011001011001110001;
#10000;
	data_in <= 24'b100100110111101101010101;
#10000;
	data_in <= 24'b100101110111111101011001;
#10000;
	data_in <= 24'b100110111000010001011110;
#10000;
	data_in <= 24'b101000001000011101100010;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101010101001001001101110;
#10000;
	data_in <= 24'b101011011001011101110001;
#10000;
	data_in <= 24'b100101000111101101010111;
#10000;
	data_in <= 24'b100110000111111101011010;
#10000;
	data_in <= 24'b100110111000001101011111;
#10000;
	data_in <= 24'b101000001000011101100010;
#10000;
	data_in <= 24'b101001001000101101100111;
#10000;
	data_in <= 24'b101001111000111001101010;
#10000;
	data_in <= 24'b101010101001001001101110;
#10000;
	data_in <= 24'b101011101001011101110011;
#10000;
	data_in <= 24'b100100110111110001010110;
#10000;
	data_in <= 24'b100101111000000001011010;
#10000;
	data_in <= 24'b100110111000010001011111;
#10000;
	data_in <= 24'b101000001000100001100010;
#10000;
	data_in <= 24'b101001001000110001100110;
#10000;
	data_in <= 24'b101001111000111001101010;
#10000;
	data_in <= 24'b101010101001001001101110;
#10000;
	data_in <= 24'b101011011001011101110011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b101100101001101101110100;
#10000;
	data_in <= 24'b101101011001111001111001;
#10000;
	data_in <= 24'b101110001010000001111101;
#10000;
	data_in <= 24'b101110101010001101111111;
#10000;
	data_in <= 24'b101111101010011010000001;
#10000;
	data_in <= 24'b110000011010100110000101;
#10000;
	data_in <= 24'b110000111010110010001000;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b101100101001101001110110;
#10000;
	data_in <= 24'b101101011001111001111001;
#10000;
	data_in <= 24'b101110001010000101111101;
#10000;
	data_in <= 24'b101110111010010010000000;
#10000;
	data_in <= 24'b101111111010011110000010;
#10000;
	data_in <= 24'b110000011010101010000110;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b101100001001100001110100;
#10000;
	data_in <= 24'b101100101001101101110111;
#10000;
	data_in <= 24'b101101101001111101111010;
#10000;
	data_in <= 24'b101110001010000101111110;
#10000;
	data_in <= 24'b101110111010010010000000;
#10000;
	data_in <= 24'b101111111010011110000011;
#10000;
	data_in <= 24'b110000101010101110000111;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b101100001001100001110100;
#10000;
	data_in <= 24'b101100101001101101110111;
#10000;
	data_in <= 24'b101101101001111101111011;
#10000;
	data_in <= 24'b101110011010001001111111;
#10000;
	data_in <= 24'b101111001010010110000010;
#10000;
	data_in <= 24'b110000001010100010000100;
#10000;
	data_in <= 24'b110000101010101110001000;
#10000;
	data_in <= 24'b110001001010110110001010;
#10000;
	data_in <= 24'b101100001001100101110101;
#10000;
	data_in <= 24'b101100111001110001111000;
#10000;
	data_in <= 24'b101101101010000001111100;
#10000;
	data_in <= 24'b101110011010001101111111;
#10000;
	data_in <= 24'b101111001010011010000010;
#10000;
	data_in <= 24'b110000001010100110000101;
#10000;
	data_in <= 24'b110000101010101110001001;
#10000;
	data_in <= 24'b110001001010111010001011;
#10000;
	data_in <= 24'b101100011001101001110101;
#10000;
	data_in <= 24'b101100111001110001111001;
#10000;
	data_in <= 24'b101101101010000001111100;
#10000;
	data_in <= 24'b101110011010001101111111;
#10000;
	data_in <= 24'b101110111010011010000011;
#10000;
	data_in <= 24'b110000001010100110000110;
#10000;
	data_in <= 24'b110000101010101110001001;
#10000;
	data_in <= 24'b110001001010111010001011;
#10000;
	data_in <= 24'b101100011001101001110110;
#10000;
	data_in <= 24'b101100111001110001111001;
#10000;
	data_in <= 24'b101101101001111101111101;
#10000;
	data_in <= 24'b101110011010001110000000;
#10000;
	data_in <= 24'b101110111010010110000011;
#10000;
	data_in <= 24'b110000001010100110000111;
#10000;
	data_in <= 24'b110000111010110010001010;
#10000;
	data_in <= 24'b110001001010111010001100;
#10000;
	data_in <= 24'b101100011001101001110110;
#10000;
	data_in <= 24'b101100111001110101111001;
#10000;
	data_in <= 24'b101101101010000001111101;
#10000;
	data_in <= 24'b101110011010001110000000;
#10000;
	data_in <= 24'b101111001010011010000100;
#10000;
	data_in <= 24'b110000001010101010000111;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110001001010111110001011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001011010111010001010;
#10000;
	data_in <= 24'b110001101011000010001101;
#10000;
	data_in <= 24'b110010011011001010001111;
#10000;
	data_in <= 24'b110010111011010110010010;
#10000;
	data_in <= 24'b110011001011011110010101;
#10000;
	data_in <= 24'b110011011011100010010111;
#10000;
	data_in <= 24'b110100001011101010011000;
#10000;
	data_in <= 24'b110100101011101110011001;
#10000;
	data_in <= 24'b110001011010111010001100;
#10000;
	data_in <= 24'b110001111011000010001111;
#10000;
	data_in <= 24'b110010101011001010010001;
#10000;
	data_in <= 24'b110011001011011010010011;
#10000;
	data_in <= 24'b110011011011100010010101;
#10000;
	data_in <= 24'b110011101011100110011000;
#10000;
	data_in <= 24'b110100001011101010011001;
#10000;
	data_in <= 24'b110100101011110010011011;
#10000;
	data_in <= 24'b110001101010111010001101;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110010101011001110010010;
#10000;
	data_in <= 24'b110010111011010110010011;
#10000;
	data_in <= 24'b110011011011100110010110;
#10000;
	data_in <= 24'b110011111011101010011001;
#10000;
	data_in <= 24'b110100011011101110011010;
#10000;
	data_in <= 24'b110100111011110110011100;
#10000;
	data_in <= 24'b110001101010111110001101;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110010101011010010010010;
#10000;
	data_in <= 24'b110011001011011010010100;
#10000;
	data_in <= 24'b110011101011100110010111;
#10000;
	data_in <= 24'b110011111011101010011010;
#10000;
	data_in <= 24'b110100011011110010011011;
#10000;
	data_in <= 24'b110100111011110110011100;
#10000;
	data_in <= 24'b110001101011000010001110;
#10000;
	data_in <= 24'b110010011011001110010001;
#10000;
	data_in <= 24'b110010101011011010010100;
#10000;
	data_in <= 24'b110011011011100010010101;
#10000;
	data_in <= 24'b110011101011100110011000;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110100011011110010011011;
#10000;
	data_in <= 24'b110100111011111010011101;
#10000;
	data_in <= 24'b110001101011000110001110;
#10000;
	data_in <= 24'b110010011011001110010001;
#10000;
	data_in <= 24'b110010101011010110010011;
#10000;
	data_in <= 24'b110011011011100010010110;
#10000;
	data_in <= 24'b110011101011100110011000;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110100101011110110011100;
#10000;
	data_in <= 24'b110101001011111110011110;
#10000;
	data_in <= 24'b110001111011000010001111;
#10000;
	data_in <= 24'b110010011011001010010010;
#10000;
	data_in <= 24'b110010101011010110010100;
#10000;
	data_in <= 24'b110011011011011110010110;
#10000;
	data_in <= 24'b110011101011100110011001;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110100101011110110011100;
#10000;
	data_in <= 24'b110101001011111110011111;
#10000;
	data_in <= 24'b110001101011000110001111;
#10000;
	data_in <= 24'b110010011011001110010010;
#10000;
	data_in <= 24'b110010101011011010010100;
#10000;
	data_in <= 24'b110011011011100010010111;
#10000;
	data_in <= 24'b110011101011100110011001;
#10000;
	data_in <= 24'b110011111011110010011010;
#10000;
	data_in <= 24'b110100101011110110011100;
#10000;
	data_in <= 24'b110101001011111110011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110100111011110110011100;
#10000;
	data_in <= 24'b110101001011111110011110;
#10000;
	data_in <= 24'b110101101100000110011111;
#10000;
	data_in <= 24'b110101111100001010100000;
#10000;
	data_in <= 24'b110110001100001110100010;
#10000;
	data_in <= 24'b110110001100001110100011;
#10000;
	data_in <= 24'b110110001100010010100100;
#10000;
	data_in <= 24'b110111001100010110100011;
#10000;
	data_in <= 24'b110101001011111010011101;
#10000;
	data_in <= 24'b110101001011111110011111;
#10000;
	data_in <= 24'b110101111100001010100000;
#10000;
	data_in <= 24'b110110001100001110100001;
#10000;
	data_in <= 24'b110110001100001110100010;
#10000;
	data_in <= 24'b110110011100010010100100;
#10000;
	data_in <= 24'b110110011100010110100101;
#10000;
	data_in <= 24'b110111001100011010100011;
#10000;
	data_in <= 24'b110101001011111010011111;
#10000;
	data_in <= 24'b110101011100000010100000;
#10000;
	data_in <= 24'b110101111100001010100001;
#10000;
	data_in <= 24'b110110001100001110100010;
#10000;
	data_in <= 24'b110110011100001110100011;
#10000;
	data_in <= 24'b110110011100010010100100;
#10000;
	data_in <= 24'b110110011100011010100111;
#10000;
	data_in <= 24'b110110111100010010100010;
#10000;
	data_in <= 24'b110101001011111110011110;
#10000;
	data_in <= 24'b110101101100000110100001;
#10000;
	data_in <= 24'b110101111100001010100001;
#10000;
	data_in <= 24'b110110001100001110100010;
#10000;
	data_in <= 24'b110110011100010010100100;
#10000;
	data_in <= 24'b110110101100010110100101;
#10000;
	data_in <= 24'b110110101100011110100111;
#10000;
	data_in <= 24'b110110111100010110100011;
#10000;
	data_in <= 24'b110101001100000010011111;
#10000;
	data_in <= 24'b110101011100001010100000;
#10000;
	data_in <= 24'b110110001100001110100011;
#10000;
	data_in <= 24'b110110001100010010100011;
#10000;
	data_in <= 24'b110110011100010110100100;
#10000;
	data_in <= 24'b110110101100011010100110;
#10000;
	data_in <= 24'b110110111100100010101000;
#10000;
	data_in <= 24'b110110111100010110100011;
#10000;
	data_in <= 24'b110101011100000010011111;
#10000;
	data_in <= 24'b110101011100001010100000;
#10000;
	data_in <= 24'b110110001100001110100011;
#10000;
	data_in <= 24'b110110001100001110100011;
#10000;
	data_in <= 24'b110110101100010110100101;
#10000;
	data_in <= 24'b110110101100011010100110;
#10000;
	data_in <= 24'b110110111100100010101000;
#10000;
	data_in <= 24'b110110111100011010100011;
#10000;
	data_in <= 24'b110101011100000010100000;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110101111100001110100011;
#10000;
	data_in <= 24'b110110001100001110100100;
#10000;
	data_in <= 24'b110110101100010110100110;
#10000;
	data_in <= 24'b110110101100011010100111;
#10000;
	data_in <= 24'b110110101100100010101000;
#10000;
	data_in <= 24'b110111001100011010100011;
#10000;
	data_in <= 24'b110101011100000110100000;
#10000;
	data_in <= 24'b110101011100001010100001;
#10000;
	data_in <= 24'b110101111100001110100011;
#10000;
	data_in <= 24'b110110001100010010100100;
#10000;
	data_in <= 24'b110110101100010110100110;
#10000;
	data_in <= 24'b110110101100011010100111;
#10000;
	data_in <= 24'b110110101100100010101000;
#10000;
	data_in <= 24'b110111011100100010100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110100011100001010101000;
#10000;
	data_in <= 24'b110000001100111111010101;
#10000;
	data_in <= 24'b110010011101100111100001;
#10000;
	data_in <= 24'b110011101101110111100100;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110010111100001010110000;
#10000;
	data_in <= 24'b110000011101000111011011;
#10000;
	data_in <= 24'b110010111101101011100001;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110001111100010010110111;
#10000;
	data_in <= 24'b110000101101001111011101;
#10000;
	data_in <= 24'b110010111101101011100001;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110001001100010010111011;
#10000;
	data_in <= 24'b110000101101001111011101;
#10000;
	data_in <= 24'b110010111101101011100001;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110011100011;
#10000;
	data_in <= 24'b110001111101100011011111;
#10000;
	data_in <= 24'b110101001110010011101010;
#10000;
	data_in <= 24'b110000111100010010111100;
#10000;
	data_in <= 24'b110000011101001011011100;
#10000;
	data_in <= 24'b110010011101100111100000;
#10000;
	data_in <= 24'b110010111101101111100010;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110001111101011111011110;
#10000;
	data_in <= 24'b101001111011100111000001;
#10000;
	data_in <= 24'b110010101101101011100000;
#10000;
	data_in <= 24'b110000101100001110111010;
#10000;
	data_in <= 24'b101111111101000111011010;
#10000;
	data_in <= 24'b110001111101100011011101;
#10000;
	data_in <= 24'b110010101101101011100000;
#10000;
	data_in <= 24'b110010101101101011100001;
#10000;
	data_in <= 24'b110010011101100111100000;
#10000;
	data_in <= 24'b110000111101001111011011;
#10000;
	data_in <= 24'b110010101101101111100001;
#10000;
	data_in <= 24'b110000101100000110110111;
#10000;
	data_in <= 24'b101111001100111011011000;
#10000;
	data_in <= 24'b110001011101010111011011;
#10000;
	data_in <= 24'b110001111101100011011110;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110000111100000010110001;
#10000;
	data_in <= 24'b101110011100101111010100;
#10000;
	data_in <= 24'b110000101101001111011001;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001111101100011011101;
#10000;
	data_in <= 24'b101111001100110111010100;
#10000;
	data_in <= 24'b101101001100010111001101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110100001101111111100111;
#10000;
	data_in <= 24'b110100101110000111101000;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110100011110000011101000;
#10000;
	data_in <= 24'b110100001101111111100110;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110001111101100011011110;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b110011111101111011100101;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010111101101111100010;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b101100001100001011001001;
#10000;
	data_in <= 24'b100110111010111010110110;
#10000;
	data_in <= 24'b110100011110000111101000;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b010101110110111001111001;
#10000;
	data_in <= 24'b101011011011111111000110;
#10000;
	data_in <= 24'b110101001110001111101010;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110010101101101111100010;
#10000;
	data_in <= 24'b101000111011011010111110;
#10000;
	data_in <= 24'b110001001101010111011100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110010111101101111100010;
#10000;
	data_in <= 24'b101111111101000011010110;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110010111101101111100010;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110100101110000111100111;
#10000;
	data_in <= 24'b110010111101110011100010;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b101101111100100011001111;
#10000;
	data_in <= 24'b101111101100111111010110;
#10000;
	data_in <= 24'b110010101101101011100000;
#10000;
	data_in <= 24'b110001111101100011011110;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110001111101100011011110;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010111101101111100001;
#10000;
	data_in <= 24'b110001101101011111011101;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b101001011011100010111111;
#10000;
	data_in <= 24'b110000101101001011011001;
#10000;
	data_in <= 24'b110001101101011111011101;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110101001110010011101011;
#10000;
	data_in <= 24'b110100111110001011101001;
#10000;
	data_in <= 24'b110011101101111011100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011011101110011100100;
#10000;
	data_in <= 24'b110101111110011011101101;
#10000;
	data_in <= 24'b100011111010001010101100;
#10000;
	data_in <= 24'b101010101011101111000100;
#10000;
	data_in <= 24'b110101101110010111101100;
#10000;
	data_in <= 24'b110011011101110011100100;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011011101110011100100;
#10000;
	data_in <= 24'b110100101110001011101001;
#10000;
	data_in <= 24'b101011011011111111000110;
#10000;
	data_in <= 24'b101110101100101111010011;
#10000;
	data_in <= 24'b110100101110001011101001;
#10000;
	data_in <= 24'b110100101110001011101000;
#10000;
	data_in <= 24'b110011101101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110100111110001111101010;
#10000;
	data_in <= 24'b110100111110001011101001;
#10000;
	data_in <= 24'b110001101101011111011110;
#10000;
	data_in <= 24'b101100011100001111001011;
#10000;
	data_in <= 24'b110011011101110111100011;
#10000;
	data_in <= 24'b110010111101110011100010;
#10000;
	data_in <= 24'b110010111101110011100011;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110010101101101011100001;
#10000;
	data_in <= 24'b110010111101101111100010;
#10000;
	data_in <= 24'b110001001101010011011011;
#10000;
	data_in <= 24'b101001001011011010111110;
#10000;
	data_in <= 24'b110011001101110011100011;
#10000;
	data_in <= 24'b110010111101101111100010;
#10000;
	data_in <= 24'b110000111101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110010111101101111100001;
#10000;
	data_in <= 24'b101101101100011111001111;
#10000;
	data_in <= 24'b110001111101011111011110;
#10000;
	data_in <= 24'b110100101110001011101000;
#10000;
	data_in <= 24'b110010111101101111100001;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110001111101011111011110;
#10000;
	data_in <= 24'b110001111101011111011110;
#10000;
	data_in <= 24'b110011001101110011100010;
#10000;
	data_in <= 24'b110001111101100011011110;
#10000;
	data_in <= 24'b110010101101101011100001;
#10000;
	data_in <= 24'b101110001100100111010001;
#10000;
	data_in <= 24'b101110011100101011010001;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101010111011100;
#10000;
	data_in <= 24'b101100001100001011001001;
#10000;
	data_in <= 24'b110000111101010011011010;
#10000;
	data_in <= 24'b110001101101011111011101;
#10000;
	data_in <= 24'b110000011101001011011001;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111111100110;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011011101110011100010;
#10000;
	data_in <= 24'b110001011101011111100010;
#10000;
	data_in <= 24'b110000011100011011000000;
#10000;
	data_in <= 24'b110100011011101010011000;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011111101111011100110;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011011101110011100011;
#10000;
	data_in <= 24'b110010001101100011100010;
#10000;
	data_in <= 24'b110000001100100111001001;
#10000;
	data_in <= 24'b110011101011101110011100;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011001101110011100100;
#10000;
	data_in <= 24'b110011101101110111100101;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110011011101110011100011;
#10000;
	data_in <= 24'b110010001101100111100001;
#10000;
	data_in <= 24'b101111111100110011001111;
#10000;
	data_in <= 24'b110011001011101110100000;
#10000;
	data_in <= 24'b110011101101111011100101;
#10000;
	data_in <= 24'b110101011110001111101010;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110010111101101111100010;
#10000;
	data_in <= 24'b110001111101100011100000;
#10000;
	data_in <= 24'b101111101100110011010001;
#10000;
	data_in <= 24'b110010101011110010100001;
#10000;
	data_in <= 24'b110010011101101011100000;
#10000;
	data_in <= 24'b101000011011010010111100;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110011011101110111100100;
#10000;
	data_in <= 24'b110010101101101011100001;
#10000;
	data_in <= 24'b110001101101011111011111;
#10000;
	data_in <= 24'b101111011100101011010001;
#10000;
	data_in <= 24'b110010011011110010100001;
#10000;
	data_in <= 24'b110001111101100011011110;
#10000;
	data_in <= 24'b101010011011101111000011;
#10000;
	data_in <= 24'b110001111101100011011111;
#10000;
	data_in <= 24'b110010101101101111100001;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110001001101010111011101;
#10000;
	data_in <= 24'b101110111100100011001101;
#10000;
	data_in <= 24'b110010101011101110100000;
#10000;
	data_in <= 24'b110010111101101111100001;
#10000;
	data_in <= 24'b110011001101110111100010;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110010001101100011011111;
#10000;
	data_in <= 24'b110001101101011011011100;
#10000;
	data_in <= 24'b110000101101001111011100;
#10000;
	data_in <= 24'b101110011100010111001000;
#10000;
	data_in <= 24'b110011001011101110011110;
#10000;
	data_in <= 24'b110001101101011111011101;
#10000;
	data_in <= 24'b110010001101100011011110;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b110001001101010011011010;
#10000;
	data_in <= 24'b101111101101000011011001;
#10000;
	data_in <= 24'b101110001100000110111111;
#10000;
	data_in <= 24'b110011101011110010011101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110100101011101110011010;
#10000;
	data_in <= 24'b110100001011101010011000;
#10000;
	data_in <= 24'b110011011011100010010111;
#10000;
	data_in <= 24'b110011001011011110010101;
#10000;
	data_in <= 24'b110010111011010110010010;
#10000;
	data_in <= 24'b110010011011001010001111;
#10000;
	data_in <= 24'b110001101011000010001101;
#10000;
	data_in <= 24'b110001011010111010001010;
#10000;
	data_in <= 24'b110100111011110010011011;
#10000;
	data_in <= 24'b110100001011101110011001;
#10000;
	data_in <= 24'b110011101011100110011000;
#10000;
	data_in <= 24'b110011011011100010010101;
#10000;
	data_in <= 24'b110011001011011010010011;
#10000;
	data_in <= 24'b110010101011001010010001;
#10000;
	data_in <= 24'b110001111011000010001111;
#10000;
	data_in <= 24'b110001011010111010001100;
#10000;
	data_in <= 24'b110101001011110110011010;
#10000;
	data_in <= 24'b110100011011101110011011;
#10000;
	data_in <= 24'b110011111011101010011001;
#10000;
	data_in <= 24'b110011011011100110010110;
#10000;
	data_in <= 24'b110010111011010110010011;
#10000;
	data_in <= 24'b110010101011001110010010;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110001101010111010001101;
#10000;
	data_in <= 24'b110101011011110110011011;
#10000;
	data_in <= 24'b110100011011110010011011;
#10000;
	data_in <= 24'b110011111011101010011010;
#10000;
	data_in <= 24'b110011101011100110010111;
#10000;
	data_in <= 24'b110011001011011010010100;
#10000;
	data_in <= 24'b110010101011010010010010;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110001101010111110001101;
#10000;
	data_in <= 24'b110101011011111010011100;
#10000;
	data_in <= 24'b110100011011110110011100;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110011101011100110011000;
#10000;
	data_in <= 24'b110011011011100010010101;
#10000;
	data_in <= 24'b110010101011011010010100;
#10000;
	data_in <= 24'b110010011011001110010001;
#10000;
	data_in <= 24'b110001101011000010001110;
#10000;
	data_in <= 24'b110101011011111110011100;
#10000;
	data_in <= 24'b110100101011110110011100;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110011101011100110011000;
#10000;
	data_in <= 24'b110011011011100010010110;
#10000;
	data_in <= 24'b110010101011010110010011;
#10000;
	data_in <= 24'b110010011011001110010001;
#10000;
	data_in <= 24'b110001101011000110001110;
#10000;
	data_in <= 24'b110101011011111110011110;
#10000;
	data_in <= 24'b110100101011110110011100;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110011101011100110011001;
#10000;
	data_in <= 24'b110011011011011110010110;
#10000;
	data_in <= 24'b110010101011010110010100;
#10000;
	data_in <= 24'b110010011011001010010010;
#10000;
	data_in <= 24'b110001111011000010001111;
#10000;
	data_in <= 24'b110101011100000010011111;
#10000;
	data_in <= 24'b110100101011110110011100;
#10000;
	data_in <= 24'b110011111011110010011010;
#10000;
	data_in <= 24'b110011101011100110011001;
#10000;
	data_in <= 24'b110011011011100010010111;
#10000;
	data_in <= 24'b110010101011011010010100;
#10000;
	data_in <= 24'b110010011011001110010010;
#10000;
	data_in <= 24'b110001101011000110001111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110000111010110010001000;
#10000;
	data_in <= 24'b110000011010100110000101;
#10000;
	data_in <= 24'b101111101010011010000001;
#10000;
	data_in <= 24'b101110101010001101111111;
#10000;
	data_in <= 24'b101110001010000001111101;
#10000;
	data_in <= 24'b101101011001111001111001;
#10000;
	data_in <= 24'b101100101001101101110100;
#10000;
	data_in <= 24'b101011111001011101110010;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110000011010101010000110;
#10000;
	data_in <= 24'b101111111010011110000010;
#10000;
	data_in <= 24'b101110111010010010000000;
#10000;
	data_in <= 24'b101110001010000101111101;
#10000;
	data_in <= 24'b101101011001111001111001;
#10000;
	data_in <= 24'b101100101001101001110110;
#10000;
	data_in <= 24'b101100001001100001110011;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110000101010101110000111;
#10000;
	data_in <= 24'b101111111010011110000011;
#10000;
	data_in <= 24'b101110111010010010000000;
#10000;
	data_in <= 24'b101110001010000101111110;
#10000;
	data_in <= 24'b101101101001111101111010;
#10000;
	data_in <= 24'b101100101001101101110111;
#10000;
	data_in <= 24'b101100001001100001110100;
#10000;
	data_in <= 24'b110001001010110110001010;
#10000;
	data_in <= 24'b110000101010101110001000;
#10000;
	data_in <= 24'b110000001010100010000100;
#10000;
	data_in <= 24'b101111001010010110000010;
#10000;
	data_in <= 24'b101110011010001001111111;
#10000;
	data_in <= 24'b101101101001111101111011;
#10000;
	data_in <= 24'b101100101001101101110111;
#10000;
	data_in <= 24'b101100001001100001110100;
#10000;
	data_in <= 24'b110001001010111010001011;
#10000;
	data_in <= 24'b110000101010101110001001;
#10000;
	data_in <= 24'b110000001010100110000101;
#10000;
	data_in <= 24'b101111001010011010000010;
#10000;
	data_in <= 24'b101110011010001101111111;
#10000;
	data_in <= 24'b101101101010000001111100;
#10000;
	data_in <= 24'b101100111001110001111000;
#10000;
	data_in <= 24'b101100001001100101110101;
#10000;
	data_in <= 24'b110001001010111010001011;
#10000;
	data_in <= 24'b110000101010101110001001;
#10000;
	data_in <= 24'b110000001010100110000110;
#10000;
	data_in <= 24'b101110111010011010000011;
#10000;
	data_in <= 24'b101110011010001101111111;
#10000;
	data_in <= 24'b101101101010000001111100;
#10000;
	data_in <= 24'b101100111001110001111001;
#10000;
	data_in <= 24'b101100011001101001110101;
#10000;
	data_in <= 24'b110001001010111010001100;
#10000;
	data_in <= 24'b110000111010110010001010;
#10000;
	data_in <= 24'b110000001010100110000111;
#10000;
	data_in <= 24'b101110111010010110000011;
#10000;
	data_in <= 24'b101110011010001110000000;
#10000;
	data_in <= 24'b101101101001111101111101;
#10000;
	data_in <= 24'b101100111001110001111001;
#10000;
	data_in <= 24'b101100011001101001110110;
#10000;
	data_in <= 24'b110001001010111110001011;
#10000;
	data_in <= 24'b110000111010110010001001;
#10000;
	data_in <= 24'b110000001010101010000111;
#10000;
	data_in <= 24'b101111001010011010000100;
#10000;
	data_in <= 24'b101110011010001110000000;
#10000;
	data_in <= 24'b101101101010000001111101;
#10000;
	data_in <= 24'b101100111001110101111001;
#10000;
	data_in <= 24'b101100011001101001110110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101011001001001101101110;
#10000;
	data_in <= 24'b101010011001000001101010;
#10000;
	data_in <= 24'b101001101000110001100110;
#10000;
	data_in <= 24'b101000111000100101100011;
#10000;
	data_in <= 24'b100111101000010101011110;
#10000;
	data_in <= 24'b100110101000001001011001;
#10000;
	data_in <= 24'b100101100111110101010110;
#10000;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b101011011001010001101111;
#10000;
	data_in <= 24'b101010011001000001101011;
#10000;
	data_in <= 24'b101001101000110101100111;
#10000;
	data_in <= 24'b101000111000100101100100;
#10000;
	data_in <= 24'b100111111000011001011111;
#10000;
	data_in <= 24'b100110101000001001011011;
#10000;
	data_in <= 24'b100101110111111001010111;
#10000;
	data_in <= 24'b100100100111100101010010;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b101010101001000001101011;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101001001000100101100101;
#10000;
	data_in <= 24'b100111111000010101100000;
#10000;
	data_in <= 24'b100110111000001101011100;
#10000;
	data_in <= 24'b100101100111111001010111;
#10000;
	data_in <= 24'b100100110111100101010010;
#10000;
	data_in <= 24'b101011011001010101110000;
#10000;
	data_in <= 24'b101010101001000101101100;
#10000;
	data_in <= 24'b101001111000111001101000;
#10000;
	data_in <= 24'b101001001000101001100101;
#10000;
	data_in <= 24'b100111111000011001100001;
#10000;
	data_in <= 24'b100110111000001101011101;
#10000;
	data_in <= 24'b100101110111111001011000;
#10000;
	data_in <= 24'b100100110111101001010011;
#10000;
	data_in <= 24'b101011011001011001110001;
#10000;
	data_in <= 24'b101010101001001001101101;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b100111111000011101100001;
#10000;
	data_in <= 24'b100110111000010001011110;
#10000;
	data_in <= 24'b100101110111111101011000;
#10000;
	data_in <= 24'b100100110111101101010100;
#10000;
	data_in <= 24'b101011011001011101110001;
#10000;
	data_in <= 24'b101010101001001001101110;
#10000;
	data_in <= 24'b101001111000111001101001;
#10000;
	data_in <= 24'b101001001000101101100110;
#10000;
	data_in <= 24'b101000001000011101100010;
#10000;
	data_in <= 24'b100110111000010001011110;
#10000;
	data_in <= 24'b100101110111111101011001;
#10000;
	data_in <= 24'b100100110111101101010101;
#10000;
	data_in <= 24'b101011101001011101110011;
#10000;
	data_in <= 24'b101010101001001001101110;
#10000;
	data_in <= 24'b101001111000111001101010;
#10000;
	data_in <= 24'b101001001000101101100111;
#10000;
	data_in <= 24'b101000001000011101100010;
#10000;
	data_in <= 24'b100110111000001101011111;
#10000;
	data_in <= 24'b100110000111111101011010;
#10000;
	data_in <= 24'b100101000111101101010111;
#10000;
	data_in <= 24'b101011011001011101110011;
#10000;
	data_in <= 24'b101010101001001001101110;
#10000;
	data_in <= 24'b101001111000111001101010;
#10000;
	data_in <= 24'b101001001000110001100110;
#10000;
	data_in <= 24'b101000001000100001100010;
#10000;
	data_in <= 24'b100110111000010001011111;
#10000;
	data_in <= 24'b100101111000000001011010;
#10000;
	data_in <= 24'b100100110111110001010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100101000111110101010111;
#10000;
	data_in <= 24'b100110001000000101011011;
#10000;
	data_in <= 24'b100111001000010001011111;
#10000;
	data_in <= 24'b101000001000100101100011;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101001111000111101101011;
#10000;
	data_in <= 24'b101010101001001101101111;
#10000;
	data_in <= 24'b101011101001100001110010;
#10000;
	data_in <= 24'b100101100111110001010111;
#10000;
	data_in <= 24'b100110101000000101011011;
#10000;
	data_in <= 24'b100111011000010001011111;
#10000;
	data_in <= 24'b101000001000100001100011;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101010011000111101101100;
#10000;
	data_in <= 24'b101010111001001101101111;
#10000;
	data_in <= 24'b101011101001100001110010;
#10000;
	data_in <= 24'b100101010111110001011000;
#10000;
	data_in <= 24'b100110101000000001011100;
#10000;
	data_in <= 24'b100111011000010001011111;
#10000;
	data_in <= 24'b101000001000100001100100;
#10000;
	data_in <= 24'b101001011000110001101000;
#10000;
	data_in <= 24'b101010011000111001101101;
#10000;
	data_in <= 24'b101010111001001101110000;
#10000;
	data_in <= 24'b101011101001100001110100;
#10000;
	data_in <= 24'b100101010111110101011001;
#10000;
	data_in <= 24'b100110101000000101011101;
#10000;
	data_in <= 24'b100111011000010101100000;
#10000;
	data_in <= 24'b101000001000100001100100;
#10000;
	data_in <= 24'b101001001000110101101001;
#10000;
	data_in <= 24'b101010001001000101101101;
#10000;
	data_in <= 24'b101010111001010001110000;
#10000;
	data_in <= 24'b101011101001011101110011;
#10000;
	data_in <= 24'b100101010111110101011000;
#10000;
	data_in <= 24'b100110101000001001011101;
#10000;
	data_in <= 24'b100111011000010101100000;
#10000;
	data_in <= 24'b101000011000100001100100;
#10000;
	data_in <= 24'b101001001000110101101001;
#10000;
	data_in <= 24'b101001111001001001101101;
#10000;
	data_in <= 24'b101010111001010001110000;
#10000;
	data_in <= 24'b101011111001011101110100;
#10000;
	data_in <= 24'b100101010111110101011000;
#10000;
	data_in <= 24'b100110101000000101011101;
#10000;
	data_in <= 24'b100111011000010101100001;
#10000;
	data_in <= 24'b101000011000100001100101;
#10000;
	data_in <= 24'b101001001000110101101010;
#10000;
	data_in <= 24'b101001111001001001101101;
#10000;
	data_in <= 24'b101010111001010001110001;
#10000;
	data_in <= 24'b101011111001011101110110;
#10000;
	data_in <= 24'b100101010111110001011000;
#10000;
	data_in <= 24'b100110101000000101011101;
#10000;
	data_in <= 24'b100111011000010101100001;
#10000;
	data_in <= 24'b101000011000100001100110;
#10000;
	data_in <= 24'b101001001000110101101010;
#10000;
	data_in <= 24'b101001111001000101101101;
#10000;
	data_in <= 24'b101010111001010001110001;
#10000;
	data_in <= 24'b101011111001011101110110;
#10000;
	data_in <= 24'b100101010111110101011001;
#10000;
	data_in <= 24'b100110101000001001011101;
#10000;
	data_in <= 24'b100111011000011101100010;
#10000;
	data_in <= 24'b101000011000101001100111;
#10000;
	data_in <= 24'b101001001000111001101011;
#10000;
	data_in <= 24'b101001111001001001101110;
#10000;
	data_in <= 24'b101010111001010101110010;
#10000;
	data_in <= 24'b101011111001100001110111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101100011001101101110110;
#10000;
	data_in <= 24'b101100111001110101111010;
#10000;
	data_in <= 24'b101101101010000101111110;
#10000;
	data_in <= 24'b101110101010010010000001;
#10000;
	data_in <= 24'b101111001010011110000100;
#10000;
	data_in <= 24'b110000001010101010000111;
#10000;
	data_in <= 24'b110000111010110110001010;
#10000;
	data_in <= 24'b110001001010111010001100;
#10000;
	data_in <= 24'b101100101001101101110111;
#10000;
	data_in <= 24'b101101001001110101111010;
#10000;
	data_in <= 24'b101101111010000001111110;
#10000;
	data_in <= 24'b101110111010001110000001;
#10000;
	data_in <= 24'b101111011010011110000100;
#10000;
	data_in <= 24'b110000001010101010000111;
#10000;
	data_in <= 24'b110000111010110110001011;
#10000;
	data_in <= 24'b110001011010111010001101;
#10000;
	data_in <= 24'b101100101001101101111000;
#10000;
	data_in <= 24'b101101001001110101111011;
#10000;
	data_in <= 24'b101101111010000001111111;
#10000;
	data_in <= 24'b101110111010001110000001;
#10000;
	data_in <= 24'b101111011010011110000101;
#10000;
	data_in <= 24'b110000001010101010001000;
#10000;
	data_in <= 24'b110000111010110110001011;
#10000;
	data_in <= 24'b110001011010111010001101;
#10000;
	data_in <= 24'b101100101001101101111000;
#10000;
	data_in <= 24'b101101001001111001111100;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101110111010010010000010;
#10000;
	data_in <= 24'b101111011010011110000101;
#10000;
	data_in <= 24'b110000001010101110001000;
#10000;
	data_in <= 24'b110000111010110110001100;
#10000;
	data_in <= 24'b110001011010111110001101;
#10000;
	data_in <= 24'b101100101001110001111001;
#10000;
	data_in <= 24'b101101011001111001111100;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101110111010010010000010;
#10000;
	data_in <= 24'b101111011010011110000110;
#10000;
	data_in <= 24'b110000001010101110001000;
#10000;
	data_in <= 24'b110000111010111010001100;
#10000;
	data_in <= 24'b110001011011000010001110;
#10000;
	data_in <= 24'b101100101001110001111010;
#10000;
	data_in <= 24'b101101011001111001111100;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101110111010010010000011;
#10000;
	data_in <= 24'b101111011010011110000110;
#10000;
	data_in <= 24'b110000001010101010001001;
#10000;
	data_in <= 24'b110000111010111010001101;
#10000;
	data_in <= 24'b110001001010111110010000;
#10000;
	data_in <= 24'b101100101001101101111001;
#10000;
	data_in <= 24'b101101011001111001111100;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101110111010010110000011;
#10000;
	data_in <= 24'b101111011010011110000110;
#10000;
	data_in <= 24'b110000001010101110001001;
#10000;
	data_in <= 24'b110000111010111010001100;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b101100101001110001111010;
#10000;
	data_in <= 24'b101101011001111101111100;
#10000;
	data_in <= 24'b101110001010001110000001;
#10000;
	data_in <= 24'b101110111010011010000100;
#10000;
	data_in <= 24'b101111011010100010000110;
#10000;
	data_in <= 24'b110000001010101110001010;
#10000;
	data_in <= 24'b110000111010110110001101;
#10000;
	data_in <= 24'b110001001011000110001111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001111011000110010000;
#10000;
	data_in <= 24'b110010011011010010010010;
#10000;
	data_in <= 24'b110010111011011010010100;
#10000;
	data_in <= 24'b110011011011100110010110;
#10000;
	data_in <= 24'b110011101011101010011001;
#10000;
	data_in <= 24'b110100001011110010011011;
#10000;
	data_in <= 24'b110100101011111010011101;
#10000;
	data_in <= 24'b110101001100000010100000;
#10000;
	data_in <= 24'b110001111011000110010000;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110010111011011010010100;
#10000;
	data_in <= 24'b110011011011100110010110;
#10000;
	data_in <= 24'b110100001011101010011001;
#10000;
	data_in <= 24'b110100011011101110011011;
#10000;
	data_in <= 24'b110100111011111010011101;
#10000;
	data_in <= 24'b110101011100000110100000;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110010111011011010010101;
#10000;
	data_in <= 24'b110011011011100110010111;
#10000;
	data_in <= 24'b110100001011101010011010;
#10000;
	data_in <= 24'b110100011011101110011100;
#10000;
	data_in <= 24'b110100111011111010011101;
#10000;
	data_in <= 24'b110101011100000110100000;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110010111011011110010101;
#10000;
	data_in <= 24'b110011011011100110010111;
#10000;
	data_in <= 24'b110100001011101110011010;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100111011111010011110;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110001111011000110010000;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110010111011100010010110;
#10000;
	data_in <= 24'b110011011011101010011000;
#10000;
	data_in <= 24'b110100001011101110011010;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100111011111010011110;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110001111011000110010010;
#10000;
	data_in <= 24'b110010101011010010010100;
#10000;
	data_in <= 24'b110010111011011110010110;
#10000;
	data_in <= 24'b110011101011100110011010;
#10000;
	data_in <= 24'b110100001011101110011011;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100111011111110011110;
#10000;
	data_in <= 24'b110101011100000110100010;
#10000;
	data_in <= 24'b110001111011000110010010;
#10000;
	data_in <= 24'b110010101011010010010100;
#10000;
	data_in <= 24'b110010111011011010010110;
#10000;
	data_in <= 24'b110011101011100110011001;
#10000;
	data_in <= 24'b110100001011101110011011;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100111011111110011111;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110001111011010010010010;
#10000;
	data_in <= 24'b110010101011010110010101;
#10000;
	data_in <= 24'b110010111011011110010111;
#10000;
	data_in <= 24'b110011101011101010011010;
#10000;
	data_in <= 24'b110100001011101110011100;
#10000;
	data_in <= 24'b110100011011110110011101;
#10000;
	data_in <= 24'b110100111100000010100000;
#10000;
	data_in <= 24'b110101011100001010100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101011100001010100010;
#10000;
	data_in <= 24'b110101011100001110100010;
#10000;
	data_in <= 24'b110101111100010010100100;
#10000;
	data_in <= 24'b110110001100010010100100;
#10000;
	data_in <= 24'b110110101100011010100110;
#10000;
	data_in <= 24'b110110101100011110101000;
#10000;
	data_in <= 24'b110110101100100010101000;
#10000;
	data_in <= 24'b110111101100100110101000;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110110001100010010100100;
#10000;
	data_in <= 24'b110110001100010010100100;
#10000;
	data_in <= 24'b110110101100010110100110;
#10000;
	data_in <= 24'b110110101100011110101000;
#10000;
	data_in <= 24'b110110101100100010101000;
#10000;
	data_in <= 24'b110111101100101010101001;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110110001100010010100100;
#10000;
	data_in <= 24'b110110001100010010100110;
#10000;
	data_in <= 24'b110110101100010110100111;
#10000;
	data_in <= 24'b110110101100011010100111;
#10000;
	data_in <= 24'b110110101100100010101001;
#10000;
	data_in <= 24'b110111101100101110101011;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110101101100001110100010;
#10000;
	data_in <= 24'b110110001100010110100101;
#10000;
	data_in <= 24'b110110001100010110100110;
#10000;
	data_in <= 24'b110110101100011010101000;
#10000;
	data_in <= 24'b110110101100011110101000;
#10000;
	data_in <= 24'b110110101100100010101001;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110101101100010010100011;
#10000;
	data_in <= 24'b110110001100010110100100;
#10000;
	data_in <= 24'b110110001100010110100110;
#10000;
	data_in <= 24'b110110101100011110101000;
#10000;
	data_in <= 24'b110110101100011110101000;
#10000;
	data_in <= 24'b110110101100100010101001;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110110001100010110100101;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110101100011110101001;
#10000;
	data_in <= 24'b110110101100011110101001;
#10000;
	data_in <= 24'b110110101100100010101010;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110110001100010110100101;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110101100011110101001;
#10000;
	data_in <= 24'b110110101100100010101001;
#10000;
	data_in <= 24'b110110101100100010101001;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110101100011010101001;
#10000;
	data_in <= 24'b110110101100100110101001;
#10000;
	data_in <= 24'b110110111100100110101010;
#10000;
	data_in <= 24'b110111001100101010101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001011011111110101100;
#10000;
	data_in <= 24'b101101011100011111001111;
#10000;
	data_in <= 24'b101111111100111111010110;
#10000;
	data_in <= 24'b110000101101001011011001;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110001011101011011011101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101010011011101111000011;
#10000;
	data_in <= 24'b110010111011111110100111;
#10000;
	data_in <= 24'b101100011100000111001000;
#10000;
	data_in <= 24'b101110111100110011010011;
#10000;
	data_in <= 24'b101111101101000011010110;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000011101001011011001;
#10000;
	data_in <= 24'b110000101101001111011001;
#10000;
	data_in <= 24'b110101001100001010100101;
#10000;
	data_in <= 24'b101100001011101110111100;
#10000;
	data_in <= 24'b101101001100011111001111;
#10000;
	data_in <= 24'b101110101100110011010010;
#10000;
	data_in <= 24'b101111001100110111010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111001100110111010011;
#10000;
	data_in <= 24'b110110111100011110100111;
#10000;
	data_in <= 24'b101101111011100010101111;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101101101100011111001101;
#10000;
	data_in <= 24'b101110001100100111010000;
#10000;
	data_in <= 24'b101110011100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110011100101011010001;
#10000;
	data_in <= 24'b110111111100101010101011;
#10000;
	data_in <= 24'b110001101011110010100101;
#10000;
	data_in <= 24'b101001101011011110111101;
#10000;
	data_in <= 24'b101100001100001011001001;
#10000;
	data_in <= 24'b101101001100010111001011;
#10000;
	data_in <= 24'b101101001100011011001101;
#10000;
	data_in <= 24'b101101011100011111001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110110011100010110100110;
#10000;
	data_in <= 24'b101011011011001010101011;
#10000;
	data_in <= 24'b101001001011100111000011;
#10000;
	data_in <= 24'b101011101100000011000110;
#10000;
	data_in <= 24'b101100001100001011001000;
#10000;
	data_in <= 24'b101100011100001111001001;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b110110111100100110101011;
#10000;
	data_in <= 24'b110111111100110010101100;
#10000;
	data_in <= 24'b110010101011110010100010;
#10000;
	data_in <= 24'b101000001010110110101111;
#10000;
	data_in <= 24'b101000111011011111000001;
#10000;
	data_in <= 24'b101010101011110011000010;
#10000;
	data_in <= 24'b101010111011110111000101;
#10000;
	data_in <= 24'b101011001011111111000110;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110111111100101110101100;
#10000;
	data_in <= 24'b110000011011011110100001;
#10000;
	data_in <= 24'b100111001010101010101101;
#10000;
	data_in <= 24'b100111011011001010111100;
#10000;
	data_in <= 24'b101001001011011110111111;
#10000;
	data_in <= 24'b101001011011100010111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001011101011011011101;
#10000;
	data_in <= 24'b110000111101010011011010;
#10000;
	data_in <= 24'b110001111101011111011110;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b100011001010000110101001;
#10000;
	data_in <= 24'b101111011100110111010100;
#10000;
	data_in <= 24'b110001001101010111011100;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000011101001111011001;
#10000;
	data_in <= 24'b101101001100010111001101;
#10000;
	data_in <= 24'b101011111100000111001000;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000111101010011011011;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b110000001101000011010111;
#10000;
	data_in <= 24'b101010111011110111000100;
#10000;
	data_in <= 24'b101000111011011110111110;
#10000;
	data_in <= 24'b110000011101001011011000;
#10000;
	data_in <= 24'b101111001100110111010011;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100110111010100;
#10000;
	data_in <= 24'b101110001100101011010000;
#10000;
	data_in <= 24'b101110111100110111010100;
#10000;
	data_in <= 24'b101111011100111011010101;
#10000;
	data_in <= 24'b101110001100101011010000;
#10000;
	data_in <= 24'b101110011100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101101011100011111001101;
#10000;
	data_in <= 24'b101101001100011011001101;
#10000;
	data_in <= 24'b101101001100011011001101;
#10000;
	data_in <= 24'b101101011100011111001110;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101011011011111111000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011011111111000111;
#10000;
	data_in <= 24'b101001111011101011000001;
#10000;
	data_in <= 24'b101001111011101011000001;
#10000;
	data_in <= 24'b101010001011101111000010;
#10000;
	data_in <= 24'b101010001011101111000010;
#10000;
	data_in <= 24'b101010001011101111000010;
#10000;
	data_in <= 24'b101010001011101111000010;
#10000;
	data_in <= 24'b101001111011101111000001;
#10000;
	data_in <= 24'b101001111011101011000001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b101111011100110111010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100110111010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110011100101011010001;
#10000;
	data_in <= 24'b101110001100101011010000;
#10000;
	data_in <= 24'b101110001100101011010000;
#10000;
	data_in <= 24'b101110011100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101101011100011111001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101001100010111001100;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101001100010111001100;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011111001110;
#10000;
	data_in <= 24'b101100011100001111001001;
#10000;
	data_in <= 24'b101100001100001011001001;
#10000;
	data_in <= 24'b101011111100000111001000;
#10000;
	data_in <= 24'b101010111011110111000101;
#10000;
	data_in <= 24'b101010111011110011000101;
#10000;
	data_in <= 24'b101100001100001011001001;
#10000;
	data_in <= 24'b101100001100001011001001;
#10000;
	data_in <= 24'b101100011100001111001010;
#10000;
	data_in <= 24'b101011001011111111000110;
#10000;
	data_in <= 24'b101010001011101111000011;
#10000;
	data_in <= 24'b101100001100001111000101;
#10000;
	data_in <= 24'b011111011000111110101101;
#10000;
	data_in <= 24'b011101001000011010101001;
#10000;
	data_in <= 24'b101100111100011011000110;
#10000;
	data_in <= 24'b101001101011100111000010;
#10000;
	data_in <= 24'b101010111011111011000101;
#10000;
	data_in <= 24'b101001001011011110111111;
#10000;
	data_in <= 24'b101010001011101110111110;
#10000;
	data_in <= 24'b101000101011010110111000;
#10000;
	data_in <= 24'b001011000011111110010000;
#10000;
	data_in <= 24'b000111110011001010001100;
#10000;
	data_in <= 24'b100110011010101110110101;
#10000;
	data_in <= 24'b101010101011110110111110;
#10000;
	data_in <= 24'b101001001011011110111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b101101001100011011001101;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110001011101011011011100;
#10000;
	data_in <= 24'b101101001100011011001100;
#10000;
	data_in <= 24'b101111101100111011010101;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b101111011100111011010101;
#10000;
	data_in <= 24'b101111111101000011010111;
#10000;
	data_in <= 24'b101111011100111111010101;
#10000;
	data_in <= 24'b110000001101000111011000;
#10000;
	data_in <= 24'b101111011100110111010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101111011100111011010101;
#10000;
	data_in <= 24'b101001011011100011000000;
#10000;
	data_in <= 24'b101100111100010111001100;
#10000;
	data_in <= 24'b110000001101000011010111;
#10000;
	data_in <= 24'b101111001100110111010011;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101110011100101111010001;
#10000;
	data_in <= 24'b101101101100100011001111;
#10000;
	data_in <= 24'b101101111100100111010000;
#10000;
	data_in <= 24'b101110011100101111010001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101101100100011001111;
#10000;
	data_in <= 24'b101101011100011111001110;
#10000;
	data_in <= 24'b101101011100011011001101;
#10000;
	data_in <= 24'b101101011100011111001101;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100011100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100101100001111001010;
#10000;
	data_in <= 24'b101100011100001111001010;
#10000;
	data_in <= 24'b101011001011111111000110;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011100000011000111;
#10000;
	data_in <= 24'b101011011011111111000110;
#10000;
	data_in <= 24'b101010111011111011000101;
#10000;
	data_in <= 24'b101001111011101011000000;
#10000;
	data_in <= 24'b101001111011101111000001;
#10000;
	data_in <= 24'b101010001011101111000010;
#10000;
	data_in <= 24'b101010001011101111000010;
#10000;
	data_in <= 24'b101001111011101111000010;
#10000;
	data_in <= 24'b101001111011101011000001;
#10000;
	data_in <= 24'b101001101011100111000000;
#10000;
	data_in <= 24'b101001011011100110111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b101100111100010011001100;
#10000;
	data_in <= 24'b110000101101001011011001;
#10000;
	data_in <= 24'b110000101101001111011010;
#10000;
	data_in <= 24'b110000001101000011010110;
#10000;
	data_in <= 24'b101110001100101111010101;
#10000;
	data_in <= 24'b101110001011110010110110;
#10000;
	data_in <= 24'b110100101011111010011101;
#10000;
	data_in <= 24'b101110111100110111010011;
#10000;
	data_in <= 24'b100011001010000010101010;
#10000;
	data_in <= 24'b101111011100110111010100;
#10000;
	data_in <= 24'b110000001101000111010111;
#10000;
	data_in <= 24'b101111001100110111010011;
#10000;
	data_in <= 24'b101100101100010111001110;
#10000;
	data_in <= 24'b101111011011100010101010;
#10000;
	data_in <= 24'b110101111100000010011110;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b110000011101001011011001;
#10000;
	data_in <= 24'b101111011100111011010100;
#10000;
	data_in <= 24'b101110111100110011010010;
#10000;
	data_in <= 24'b101101101100100111010000;
#10000;
	data_in <= 24'b101011011011110111000001;
#10000;
	data_in <= 24'b110001101011100010011111;
#10000;
	data_in <= 24'b110110001100001110100001;
#10000;
	data_in <= 24'b101110001100101011010001;
#10000;
	data_in <= 24'b101101111100100111001111;
#10000;
	data_in <= 24'b101101111100100111010000;
#10000;
	data_in <= 24'b101101011100011111001101;
#10000;
	data_in <= 24'b101011101100001011001010;
#10000;
	data_in <= 24'b101100001011010110101110;
#10000;
	data_in <= 24'b110100101011111110011101;
#10000;
	data_in <= 24'b110101111100010010100011;
#10000;
	data_in <= 24'b101101011100011111001101;
#10000;
	data_in <= 24'b101101001100011011001101;
#10000;
	data_in <= 24'b101100111100010011001011;
#10000;
	data_in <= 24'b101011111100000111001001;
#10000;
	data_in <= 24'b101001011011011010111100;
#10000;
	data_in <= 24'b110000011011011010011101;
#10000;
	data_in <= 24'b110110011100010110100011;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b101100011100001011001001;
#10000;
	data_in <= 24'b101011111100000111001000;
#10000;
	data_in <= 24'b101011011011111111000110;
#10000;
	data_in <= 24'b101000111011011011000000;
#10000;
	data_in <= 24'b101100001011000010100011;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b101010101011110111000011;
#10000;
	data_in <= 24'b101010011011101011000010;
#10000;
	data_in <= 24'b101000001011010010111110;
#10000;
	data_in <= 24'b101001101010110010100101;
#10000;
	data_in <= 24'b110011101011110110011110;
#10000;
	data_in <= 24'b110110011100011010100111;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b101001001011011110111111;
#10000;
	data_in <= 24'b100110101010111010110111;
#10000;
	data_in <= 24'b101001011010101010100010;
#10000;
	data_in <= 24'b110011001011101110011110;
#10000;
	data_in <= 24'b110110111100011110101001;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101011100001010100001;
#10000;
	data_in <= 24'b110100101011111010011101;
#10000;
	data_in <= 24'b110100001011110010011011;
#10000;
	data_in <= 24'b110011101011101010011001;
#10000;
	data_in <= 24'b110011011011100110010110;
#10000;
	data_in <= 24'b110010111011011010010100;
#10000;
	data_in <= 24'b110010011011010010010010;
#10000;
	data_in <= 24'b110001111011000110010000;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110100111011111010011101;
#10000;
	data_in <= 24'b110100011011101110011011;
#10000;
	data_in <= 24'b110100001011101010011001;
#10000;
	data_in <= 24'b110011011011100110010110;
#10000;
	data_in <= 24'b110010111011011010010100;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110001111011000110010000;
#10000;
	data_in <= 24'b110101001100000110100001;
#10000;
	data_in <= 24'b110100111011111010011101;
#10000;
	data_in <= 24'b110100011011101110011100;
#10000;
	data_in <= 24'b110100001011101010011010;
#10000;
	data_in <= 24'b110011011011100110010111;
#10000;
	data_in <= 24'b110010111011011010010101;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110101011100000010100001;
#10000;
	data_in <= 24'b110100111011111010011110;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100001011101110011010;
#10000;
	data_in <= 24'b110011011011100110010111;
#10000;
	data_in <= 24'b110010111011011110010101;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110010001011000110010000;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110100111011111010011110;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100001011101110011010;
#10000;
	data_in <= 24'b110011011011101010011000;
#10000;
	data_in <= 24'b110010111011100010010110;
#10000;
	data_in <= 24'b110010101011010010010011;
#10000;
	data_in <= 24'b110001111011000110010000;
#10000;
	data_in <= 24'b110101011100000110100010;
#10000;
	data_in <= 24'b110100111011111110011110;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100001011101110011011;
#10000;
	data_in <= 24'b110011101011100110011010;
#10000;
	data_in <= 24'b110010111011011110010110;
#10000;
	data_in <= 24'b110010101011010010010100;
#10000;
	data_in <= 24'b110001111011000110010010;
#10000;
	data_in <= 24'b110101011100000110100001;
#10000;
	data_in <= 24'b110100111011111110011111;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100001011101110011011;
#10000;
	data_in <= 24'b110011101011100110011001;
#10000;
	data_in <= 24'b110010111011011010010110;
#10000;
	data_in <= 24'b110010101011010010010100;
#10000;
	data_in <= 24'b110001111011000110010010;
#10000;
	data_in <= 24'b110101011100001010100010;
#10000;
	data_in <= 24'b110100111100000010100000;
#10000;
	data_in <= 24'b110100011011110110011101;
#10000;
	data_in <= 24'b110100001011101110011100;
#10000;
	data_in <= 24'b110011101011101010011010;
#10000;
	data_in <= 24'b110010111011011110010111;
#10000;
	data_in <= 24'b110010101011010110010101;
#10000;
	data_in <= 24'b110001111011010010010010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001001010111010001100;
#10000;
	data_in <= 24'b110000111010110110001010;
#10000;
	data_in <= 24'b110000001010101010000111;
#10000;
	data_in <= 24'b101111001010011110000100;
#10000;
	data_in <= 24'b101110101010010010000001;
#10000;
	data_in <= 24'b101101101010000101111110;
#10000;
	data_in <= 24'b101100111001110101111010;
#10000;
	data_in <= 24'b101100011001101101110110;
#10000;
	data_in <= 24'b110001011010111010001101;
#10000;
	data_in <= 24'b110000111010110110001011;
#10000;
	data_in <= 24'b110000001010101010000111;
#10000;
	data_in <= 24'b101111011010011110000100;
#10000;
	data_in <= 24'b101110111010001110000001;
#10000;
	data_in <= 24'b101101111010000001111110;
#10000;
	data_in <= 24'b101101001001110101111010;
#10000;
	data_in <= 24'b101100101001101101110111;
#10000;
	data_in <= 24'b110001011010111010001101;
#10000;
	data_in <= 24'b110000111010110110001011;
#10000;
	data_in <= 24'b110000001010101010001000;
#10000;
	data_in <= 24'b101111011010011110000101;
#10000;
	data_in <= 24'b101110111010001110000001;
#10000;
	data_in <= 24'b101110001010000001111111;
#10000;
	data_in <= 24'b101101001001110101111011;
#10000;
	data_in <= 24'b101100101001101101111000;
#10000;
	data_in <= 24'b110001011010111110001101;
#10000;
	data_in <= 24'b110000111010110110001100;
#10000;
	data_in <= 24'b110000001010101110001000;
#10000;
	data_in <= 24'b101111011010011110000101;
#10000;
	data_in <= 24'b101110111010010010000010;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101101001001111001111100;
#10000;
	data_in <= 24'b101100101001101101111000;
#10000;
	data_in <= 24'b110001011011000010001110;
#10000;
	data_in <= 24'b110000111010111010001100;
#10000;
	data_in <= 24'b110000001010101110001000;
#10000;
	data_in <= 24'b101111011010011110000110;
#10000;
	data_in <= 24'b101110111010010010000010;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101101011001111001111100;
#10000;
	data_in <= 24'b101100101001110001111001;
#10000;
	data_in <= 24'b110001001010111110010000;
#10000;
	data_in <= 24'b110000111010111010001101;
#10000;
	data_in <= 24'b110000001010101010001001;
#10000;
	data_in <= 24'b101111011010011110000110;
#10000;
	data_in <= 24'b101110111010010010000011;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101101011001111001111100;
#10000;
	data_in <= 24'b101100101001110001111010;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110000111010111010001100;
#10000;
	data_in <= 24'b110000001010101110001001;
#10000;
	data_in <= 24'b101111011010011110000110;
#10000;
	data_in <= 24'b101110111010010110000011;
#10000;
	data_in <= 24'b101110001010000101111111;
#10000;
	data_in <= 24'b101101011001111001111100;
#10000;
	data_in <= 24'b101100101001101101111001;
#10000;
	data_in <= 24'b110001001011000110001111;
#10000;
	data_in <= 24'b110000111010110110001101;
#10000;
	data_in <= 24'b110000001010101110001010;
#10000;
	data_in <= 24'b101111011010100010000110;
#10000;
	data_in <= 24'b101110111010011010000100;
#10000;
	data_in <= 24'b101110001010001110000001;
#10000;
	data_in <= 24'b101101011001111101111100;
#10000;
	data_in <= 24'b101100101001110001111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101011101001100001110010;
#10000;
	data_in <= 24'b101010101001001101101111;
#10000;
	data_in <= 24'b101001111000111101101011;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101000001000100101100011;
#10000;
	data_in <= 24'b100111001000010001011111;
#10000;
	data_in <= 24'b100110001000000101011011;
#10000;
	data_in <= 24'b100101000111110101010111;
#10000;
	data_in <= 24'b101011101001100001110010;
#10000;
	data_in <= 24'b101010111001001101101111;
#10000;
	data_in <= 24'b101010011000111101101100;
#10000;
	data_in <= 24'b101001001000110001100111;
#10000;
	data_in <= 24'b101000001000100001100011;
#10000;
	data_in <= 24'b100111011000010001011111;
#10000;
	data_in <= 24'b100110101000000101011011;
#10000;
	data_in <= 24'b100101100111110001010111;
#10000;
	data_in <= 24'b101011101001100001110100;
#10000;
	data_in <= 24'b101010111001001101110000;
#10000;
	data_in <= 24'b101010011000111001101101;
#10000;
	data_in <= 24'b101001011000110001101000;
#10000;
	data_in <= 24'b101000001000100001100100;
#10000;
	data_in <= 24'b100111011000010001011111;
#10000;
	data_in <= 24'b100110101000000001011100;
#10000;
	data_in <= 24'b100101010111110001011000;
#10000;
	data_in <= 24'b101011101001011101110011;
#10000;
	data_in <= 24'b101010111001010001110000;
#10000;
	data_in <= 24'b101010001001000101101101;
#10000;
	data_in <= 24'b101001001000110101101001;
#10000;
	data_in <= 24'b101000001000100001100100;
#10000;
	data_in <= 24'b100111011000010101100000;
#10000;
	data_in <= 24'b100110101000000101011101;
#10000;
	data_in <= 24'b100101010111110101011001;
#10000;
	data_in <= 24'b101011111001011101110100;
#10000;
	data_in <= 24'b101010111001010001110000;
#10000;
	data_in <= 24'b101001111001001001101101;
#10000;
	data_in <= 24'b101001001000110101101001;
#10000;
	data_in <= 24'b101000011000100001100100;
#10000;
	data_in <= 24'b100111011000010101100000;
#10000;
	data_in <= 24'b100110101000001001011101;
#10000;
	data_in <= 24'b100101010111110101011000;
#10000;
	data_in <= 24'b101011111001011101110110;
#10000;
	data_in <= 24'b101010111001010001110001;
#10000;
	data_in <= 24'b101001111001001001101101;
#10000;
	data_in <= 24'b101001001000110101101010;
#10000;
	data_in <= 24'b101000011000100001100101;
#10000;
	data_in <= 24'b100111011000010101100001;
#10000;
	data_in <= 24'b100110101000000101011101;
#10000;
	data_in <= 24'b100101010111110101011000;
#10000;
	data_in <= 24'b101011111001011101110110;
#10000;
	data_in <= 24'b101010111001010001110001;
#10000;
	data_in <= 24'b101001111001000101101101;
#10000;
	data_in <= 24'b101001001000110101101010;
#10000;
	data_in <= 24'b101000011000100001100110;
#10000;
	data_in <= 24'b100111011000010101100001;
#10000;
	data_in <= 24'b100110101000000101011101;
#10000;
	data_in <= 24'b100101010111110001011000;
#10000;
	data_in <= 24'b101011111001100001110111;
#10000;
	data_in <= 24'b101010111001010101110010;
#10000;
	data_in <= 24'b101001111001001001101110;
#10000;
	data_in <= 24'b101001001000111001101011;
#10000;
	data_in <= 24'b101000011000101001100111;
#10000;
	data_in <= 24'b100111011000011101100010;
#10000;
	data_in <= 24'b100110101000001001011101;
#10000;
	data_in <= 24'b100101010111110101011001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100101010111110101011010;
#10000;
	data_in <= 24'b100110101000001101011110;
#10000;
	data_in <= 24'b100111011000011101100011;
#10000;
	data_in <= 24'b101000011000101101100110;
#10000;
	data_in <= 24'b101001001000111001101010;
#10000;
	data_in <= 24'b101010001001000101101110;
#10000;
	data_in <= 24'b101010111001010101110010;
#10000;
	data_in <= 24'b101011111001100101110111;
#10000;
	data_in <= 24'b100101100111110101011011;
#10000;
	data_in <= 24'b100110101000001001011111;
#10000;
	data_in <= 24'b100111011000011101100011;
#10000;
	data_in <= 24'b101000011000101001100111;
#10000;
	data_in <= 24'b101001001000111001101011;
#10000;
	data_in <= 24'b101001111001000101101111;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101011101001100001110111;
#10000;
	data_in <= 24'b100101100111111001011100;
#10000;
	data_in <= 24'b100110101000001001100000;
#10000;
	data_in <= 24'b100111101000011101100100;
#10000;
	data_in <= 24'b101000011000101101101000;
#10000;
	data_in <= 24'b101001011000111001101011;
#10000;
	data_in <= 24'b101010001001001001101111;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101100001001100101110110;
#10000;
	data_in <= 24'b100101101000000001011011;
#10000;
	data_in <= 24'b100110111000010001011111;
#10000;
	data_in <= 24'b100111101000100001100011;
#10000;
	data_in <= 24'b101000101000110001100111;
#10000;
	data_in <= 24'b101001011000111101101011;
#10000;
	data_in <= 24'b101010001001001001101111;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101100001001101001110110;
#10000;
	data_in <= 24'b100101100111111101011011;
#10000;
	data_in <= 24'b100110111000001101100000;
#10000;
	data_in <= 24'b100111101000011101100100;
#10000;
	data_in <= 24'b101000011000101101101000;
#10000;
	data_in <= 24'b101001011000111101101100;
#10000;
	data_in <= 24'b101010001001001001110000;
#10000;
	data_in <= 24'b101010111001010101110100;
#10000;
	data_in <= 24'b101100001001100101110111;
#10000;
	data_in <= 24'b100101100111111101011011;
#10000;
	data_in <= 24'b100110111000010001100000;
#10000;
	data_in <= 24'b100111101000011101100100;
#10000;
	data_in <= 24'b101000011000101101101001;
#10000;
	data_in <= 24'b101001011000111101101101;
#10000;
	data_in <= 24'b101010001001001001101111;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101011111001100101111000;
#10000;
	data_in <= 24'b100101100111111101011100;
#10000;
	data_in <= 24'b100110111000001101100001;
#10000;
	data_in <= 24'b100111101000011101100101;
#10000;
	data_in <= 24'b101000011000101101101001;
#10000;
	data_in <= 24'b101001011000111101101101;
#10000;
	data_in <= 24'b101010001001001001110001;
#10000;
	data_in <= 24'b101010111001010101110100;
#10000;
	data_in <= 24'b101011111001100101111000;
#10000;
	data_in <= 24'b100101101000000001011110;
#10000;
	data_in <= 24'b100110111000010001100010;
#10000;
	data_in <= 24'b100111101000011101100110;
#10000;
	data_in <= 24'b101000011000101101101001;
#10000;
	data_in <= 24'b101001011001000001101101;
#10000;
	data_in <= 24'b101010001001001001110010;
#10000;
	data_in <= 24'b101010111001011001110100;
#10000;
	data_in <= 24'b101100001001101001111001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101100101001110001111010;
#10000;
	data_in <= 24'b101101001010000001111100;
#10000;
	data_in <= 24'b101110001010001110000000;
#10000;
	data_in <= 24'b101110111010011010000100;
#10000;
	data_in <= 24'b101111011010100010000110;
#10000;
	data_in <= 24'b110000001010101110001010;
#10000;
	data_in <= 24'b110000111010110110001110;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b101100101001110001111011;
#10000;
	data_in <= 24'b101101011001111101111101;
#10000;
	data_in <= 24'b101110001010001110000001;
#10000;
	data_in <= 24'b101110111010011010000101;
#10000;
	data_in <= 24'b101111011010100010000111;
#10000;
	data_in <= 24'b110000001010101110001010;
#10000;
	data_in <= 24'b110000111010111010001110;
#10000;
	data_in <= 24'b110001011010111110010000;
#10000;
	data_in <= 24'b101101001001110001111011;
#10000;
	data_in <= 24'b101101101001111101111110;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101111101010100110000111;
#10000;
	data_in <= 24'b110000011010101110001010;
#10000;
	data_in <= 24'b110001001010111010001110;
#10000;
	data_in <= 24'b110001011011000010010000;
#10000;
	data_in <= 24'b101101001001110101111010;
#10000;
	data_in <= 24'b101101101010000001111110;
#10000;
	data_in <= 24'b101110011010001110000001;
#10000;
	data_in <= 24'b101111001010011010000100;
#10000;
	data_in <= 24'b101111101010100110000111;
#10000;
	data_in <= 24'b110000011010110010001011;
#10000;
	data_in <= 24'b110001001010111110001110;
#10000;
	data_in <= 24'b110001011011001010010000;
#10000;
	data_in <= 24'b101101001001111001111011;
#10000;
	data_in <= 24'b101101101010000001111110;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101111101010100110001000;
#10000;
	data_in <= 24'b110000011010110010001100;
#10000;
	data_in <= 24'b110001001011000010001110;
#10000;
	data_in <= 24'b110001011011000110010000;
#10000;
	data_in <= 24'b101101001001111001111011;
#10000;
	data_in <= 24'b101101101010000001111110;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101111101010100010001000;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110001011011000110010000;
#10000;
	data_in <= 24'b101101001001111001111100;
#10000;
	data_in <= 24'b101101101010000001111111;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101111101010100010001001;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110001011011000110010001;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b101101101010000101111111;
#10000;
	data_in <= 24'b101110011010010010000010;
#10000;
	data_in <= 24'b101111001010011010000110;
#10000;
	data_in <= 24'b101111101010100110001001;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110001011011001010010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001111011001110010010;
#10000;
	data_in <= 24'b110010011011011010010100;
#10000;
	data_in <= 24'b110010111011011110010111;
#10000;
	data_in <= 24'b110011101011101010011001;
#10000;
	data_in <= 24'b110100001011101110011100;
#10000;
	data_in <= 24'b110100011011110110011101;
#10000;
	data_in <= 24'b110100111100000010100000;
#10000;
	data_in <= 24'b110101011100001010100010;
#10000;
	data_in <= 24'b110001101011001110010010;
#10000;
	data_in <= 24'b110010011011011010010101;
#10000;
	data_in <= 24'b110010111011011110011000;
#10000;
	data_in <= 24'b110011101011101010011010;
#10000;
	data_in <= 24'b110100001011101110011100;
#10000;
	data_in <= 24'b110100011011110010011101;
#10000;
	data_in <= 24'b110100111100000010100000;
#10000;
	data_in <= 24'b110101011100001010100011;
#10000;
	data_in <= 24'b110001111011001110010010;
#10000;
	data_in <= 24'b110010101011011010010101;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110011111011101010011011;
#10000;
	data_in <= 24'b110100011011101110011100;
#10000;
	data_in <= 24'b110100101011110110011101;
#10000;
	data_in <= 24'b110101001100000010100000;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110010001011010010010011;
#10000;
	data_in <= 24'b110010101011011110010101;
#10000;
	data_in <= 24'b110011011011100110011000;
#10000;
	data_in <= 24'b110100001011101110011011;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100101011111010011110;
#10000;
	data_in <= 24'b110101001100000010100000;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110001111011001110010011;
#10000;
	data_in <= 24'b110010101011011010010110;
#10000;
	data_in <= 24'b110011001011100010011000;
#10000;
	data_in <= 24'b110011111011101110011011;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100101011111010011111;
#10000;
	data_in <= 24'b110101001100000010100001;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110001111011010010010011;
#10000;
	data_in <= 24'b110010101011011010010111;
#10000;
	data_in <= 24'b110011001011100110011000;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100101011111010011111;
#10000;
	data_in <= 24'b110101001100000010100001;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110001111011001110010100;
#10000;
	data_in <= 24'b110010101011010110010111;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110011101011101010011011;
#10000;
	data_in <= 24'b110100001011110010011101;
#10000;
	data_in <= 24'b110100101011111010011111;
#10000;
	data_in <= 24'b110101001100000010100010;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110001111011010010010100;
#10000;
	data_in <= 24'b110010101011011010010111;
#10000;
	data_in <= 24'b110011011011100010011010;
#10000;
	data_in <= 24'b110011111011101010011100;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110100101011111110011111;
#10000;
	data_in <= 24'b110101001100000110100001;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110101100011010101001;
#10000;
	data_in <= 24'b110110101100100010101001;
#10000;
	data_in <= 24'b110110111100100110101010;
#10000;
	data_in <= 24'b110111001100101010101011;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110101100011010101001;
#10000;
	data_in <= 24'b110110101100100010101010;
#10000;
	data_in <= 24'b110110111100100110101011;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110101111100001110100100;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b110110011100010110100111;
#10000;
	data_in <= 24'b110110011100010110100111;
#10000;
	data_in <= 24'b110110111100011110101001;
#10000;
	data_in <= 24'b110110111100100010101010;
#10000;
	data_in <= 24'b110111001100100010101011;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110101111100010010100100;
#10000;
	data_in <= 24'b110101111100010110100101;
#10000;
	data_in <= 24'b110110011100011010100111;
#10000;
	data_in <= 24'b110110011100011010100111;
#10000;
	data_in <= 24'b110110111100100010101000;
#10000;
	data_in <= 24'b110110111100100110101001;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110101111100001110100100;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110111100011110101001;
#10000;
	data_in <= 24'b110110111100100110101010;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110101111100001110100100;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110111100100010101010;
#10000;
	data_in <= 24'b110110111100100110101010;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110101111100001110100101;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110111100100010101001;
#10000;
	data_in <= 24'b110110111100100110101011;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110101100100010101001;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110111001100101010101011;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110111101100101110101100;
#10000;
	data_in <= 24'b110000111011100110100000;
#10000;
	data_in <= 24'b101000001010100010100011;
#10000;
	data_in <= 24'b100110011010101110110001;
#10000;
	data_in <= 24'b100111101011000110111000;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110111011100101110101111;
#10000;
	data_in <= 24'b111000001100110110101111;
#10000;
	data_in <= 24'b110100111100001010100101;
#10000;
	data_in <= 24'b100011111001101010011100;
#10000;
	data_in <= 24'b100000111001100010100011;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110111101100101110101101;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111001100101010101110;
#10000;
	data_in <= 24'b111000101100111110110000;
#10000;
	data_in <= 24'b110100001100010010101110;
#10000;
	data_in <= 24'b100011111010001010101011;
#10000;
	data_in <= 24'b100100011010010110110000;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110111101100101110101101;
#10000;
	data_in <= 24'b110111101100101110101101;
#10000;
	data_in <= 24'b110111011100101010101110;
#10000;
	data_in <= 24'b111001001101000010101111;
#10000;
	data_in <= 24'b101101111011011010101010;
#10000;
	data_in <= 24'b100010111010001010101111;
#10000;
	data_in <= 24'b100111111011001010111100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111101100101110101111;
#10000;
	data_in <= 24'b111000011100110110101111;
#10000;
	data_in <= 24'b101001111010111010101001;
#10000;
	data_in <= 24'b100011011010010010110010;
#10000;
	data_in <= 24'b101000001011001110111100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111111100110010101111;
#10000;
	data_in <= 24'b110111101100110010101110;
#10000;
	data_in <= 24'b100111111010100110101001;
#10000;
	data_in <= 24'b100011111010011010110011;
#10000;
	data_in <= 24'b101000011011010010111101;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111011100101110101111;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111011100101110101111;
#10000;
	data_in <= 24'b100111001010100010101001;
#10000;
	data_in <= 24'b100100001010011010110100;
#10000;
	data_in <= 24'b101000101011010010111101;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110111101100110010101110;
#10000;
	data_in <= 24'b110111101100101110101111;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b100111011010100010101001;
#10000;
	data_in <= 24'b100100001010011010110011;
#10000;
	data_in <= 24'b101000011011001110111101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000001011001110111010;
#10000;
	data_in <= 24'b101000011011010010111011;
#10000;
	data_in <= 24'b101000011011010010111011;
#10000;
	data_in <= 24'b101000011011010110111100;
#10000;
	data_in <= 24'b101000011011010110111100;
#10000;
	data_in <= 24'b101000011011010010111100;
#10000;
	data_in <= 24'b101000001011010010111010;
#10000;
	data_in <= 24'b100111101011000110111000;
#10000;
	data_in <= 24'b100011111010001010101001;
#10000;
	data_in <= 24'b100100011010010010101100;
#10000;
	data_in <= 24'b100100111010011110101111;
#10000;
	data_in <= 24'b100101001010100010101111;
#10000;
	data_in <= 24'b100101011010100010101111;
#10000;
	data_in <= 24'b100101001010011110101110;
#10000;
	data_in <= 24'b100100101010010110101101;
#10000;
	data_in <= 24'b100100001010010010101101;
#10000;
	data_in <= 24'b100101001010011110110000;
#10000;
	data_in <= 24'b100100101010010110101111;
#10000;
	data_in <= 24'b100100101010010110101111;
#10000;
	data_in <= 24'b100100101010011010110000;
#10000;
	data_in <= 24'b100101001010100110110010;
#10000;
	data_in <= 24'b100101111010110010110110;
#10000;
	data_in <= 24'b100111011011000110111100;
#10000;
	data_in <= 24'b101001111011110011000111;
#10000;
	data_in <= 24'b101001011011100011000010;
#10000;
	data_in <= 24'b101010001011101111000101;
#10000;
	data_in <= 24'b101010101011110111001000;
#10000;
	data_in <= 24'b101011011100000111001011;
#10000;
	data_in <= 24'b101011111100010011001110;
#10000;
	data_in <= 24'b101100111100100011010010;
#10000;
	data_in <= 24'b101101101100110011010110;
#10000;
	data_in <= 24'b101101111100111011011010;
#10000;
	data_in <= 24'b101000111011011011000000;
#10000;
	data_in <= 24'b101001101011101011000100;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101011011100001011001100;
#10000;
	data_in <= 24'b101100001100010111001111;
#10000;
	data_in <= 24'b101100111100100011010010;
#10000;
	data_in <= 24'b101101011100101111010101;
#10000;
	data_in <= 24'b101110011100110011010100;
#10000;
	data_in <= 24'b101001001011011111000001;
#10000;
	data_in <= 24'b101001111011101111000100;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101011011100000111001011;
#10000;
	data_in <= 24'b101100001100010111001111;
#10000;
	data_in <= 24'b101100111100100111010011;
#10000;
	data_in <= 24'b101110101100110011010100;
#10000;
	data_in <= 24'b110001111101001011011000;
#10000;
	data_in <= 24'b101001001011011111000001;
#10000;
	data_in <= 24'b101001111011101111000100;
#10000;
	data_in <= 24'b101010101011111011001001;
#10000;
	data_in <= 24'b101011011100000111001100;
#10000;
	data_in <= 24'b101100001100011011010000;
#10000;
	data_in <= 24'b101100111100100011010010;
#10000;
	data_in <= 24'b110000111100111111010111;
#10000;
	data_in <= 24'b110100001101101011011111;
#10000;
	data_in <= 24'b101001001011011011000001;
#10000;
	data_in <= 24'b101001111011101111000100;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101011011100001011001011;
#10000;
	data_in <= 24'b101011111100010111001111;
#10000;
	data_in <= 24'b101101001100100111010010;
#10000;
	data_in <= 24'b110010011101010011011011;
#10000;
	data_in <= 24'b110100111101110111100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100111011011000010110101;
#10000;
	data_in <= 24'b100010111001111110101110;
#10000;
	data_in <= 24'b001110100101000010011000;
#10000;
	data_in <= 24'b000001100001110110001101;
#10000;
	data_in <= 24'b000001000001110010001110;
#10000;
	data_in <= 24'b001010110100000110010101;
#10000;
	data_in <= 24'b011111111001001110101010;
#10000;
	data_in <= 24'b100111011010111110110100;
#10000;
	data_in <= 24'b100110011010110110110010;
#10000;
	data_in <= 24'b010000100101101010011101;
#10000;
	data_in <= 24'b000000000001101010010001;
#10000;
	data_in <= 24'b000100010010110010011010;
#10000;
	data_in <= 24'b000100000010110010011011;
#10000;
	data_in <= 24'b000001000001111110010100;
#10000;
	data_in <= 24'b000111100011011110010101;
#10000;
	data_in <= 24'b100010001001110110101110;
#10000;
	data_in <= 24'b101110001100111111010100;
#10000;
	data_in <= 24'b010011010110100110101101;
#10000;
	data_in <= 24'b000010000010011010011001;
#10000;
	data_in <= 24'b000101100011010010100010;
#10000;
	data_in <= 24'b000101000011001110100010;
#10000;
	data_in <= 24'b000011110010110110011101;
#10000;
	data_in <= 24'b000111110011110010011110;
#10000;
	data_in <= 24'b101000111011101011001010;
#10000;
	data_in <= 24'b110001011101100111011011;
#10000;
	data_in <= 24'b011101101000110110111000;
#10000;
	data_in <= 24'b000001110010100010011011;
#10000;
	data_in <= 24'b000100010011001010100100;
#10000;
	data_in <= 24'b000100010011001110100101;
#10000;
	data_in <= 24'b000001000010011010011101;
#10000;
	data_in <= 24'b010100010110101110101011;
#10000;
	data_in <= 24'b101111011101001011010111;
#10000;
	data_in <= 24'b110001011101000111010111;
#10000;
	data_in <= 24'b101111011100100111010000;
#10000;
	data_in <= 24'b010110000111000110101110;
#10000;
	data_in <= 24'b001000110100001110100011;
#10000;
	data_in <= 24'b001010010100100010100101;
#10000;
	data_in <= 24'b010110010111001010101101;
#10000;
	data_in <= 24'b101100111100000011001010;
#10000;
	data_in <= 24'b110000111101000111010110;
#10000;
	data_in <= 24'b110011111101100011011110;
#10000;
	data_in <= 24'b110101011101111111100010;
#10000;
	data_in <= 24'b110100001101101011011100;
#10000;
	data_in <= 24'b101110011100011011010000;
#10000;
	data_in <= 24'b101111011100100111010001;
#10000;
	data_in <= 24'b110100111101110011011101;
#10000;
	data_in <= 24'b110101011101111111100010;
#10000;
	data_in <= 24'b110011011101011111011100;
#10000;
	data_in <= 24'b110101001101111011100011;
#10000;
	data_in <= 24'b110101101110000011100101;
#10000;
	data_in <= 24'b110110011110010011101001;
#10000;
	data_in <= 24'b110111101110100111101100;
#10000;
	data_in <= 24'b110111011110100011101100;
#10000;
	data_in <= 24'b110110011110010011101001;
#10000;
	data_in <= 24'b110101101110000011100110;
#10000;
	data_in <= 24'b110101001101111011100011;
#10000;
	data_in <= 24'b110101101110000011100101;
#10000;
	data_in <= 24'b110110011110001111101000;
#10000;
	data_in <= 24'b110110111110011011101011;
#10000;
	data_in <= 24'b110111001110011111101100;
#10000;
	data_in <= 24'b110111001110011111101100;
#10000;
	data_in <= 24'b110110111110011011101011;
#10000;
	data_in <= 24'b110110001110001111101000;
#10000;
	data_in <= 24'b110101101110000011100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100111101011000010111000;
#10000;
	data_in <= 24'b101000001011001110111010;
#10000;
	data_in <= 24'b101000011011010010111011;
#10000;
	data_in <= 24'b101000011011010010111100;
#10000;
	data_in <= 24'b101000011011010010111011;
#10000;
	data_in <= 24'b101000001011010010111010;
#10000;
	data_in <= 24'b101000001011001110111001;
#10000;
	data_in <= 24'b100110101010111010110101;
#10000;
	data_in <= 24'b100101011010100110101111;
#10000;
	data_in <= 24'b100100001010010010101101;
#10000;
	data_in <= 24'b100101001010011110101110;
#10000;
	data_in <= 24'b100101001010011110101111;
#10000;
	data_in <= 24'b100101001010011110101110;
#10000;
	data_in <= 24'b100100011010010110101100;
#10000;
	data_in <= 24'b100011101010000110101001;
#10000;
	data_in <= 24'b100001101001101110100101;
#10000;
	data_in <= 24'b101011101100001111001100;
#10000;
	data_in <= 24'b100111011011001010111101;
#10000;
	data_in <= 24'b100110001010110010110110;
#10000;
	data_in <= 24'b100101001010100010110010;
#10000;
	data_in <= 24'b100100111010011010110000;
#10000;
	data_in <= 24'b100100111010011110110001;
#10000;
	data_in <= 24'b100101111010101110110101;
#10000;
	data_in <= 24'b100111001010111010111001;
#10000;
	data_in <= 24'b101110001100111011011001;
#10000;
	data_in <= 24'b101101101100101111010101;
#10000;
	data_in <= 24'b101100111100011111010010;
#10000;
	data_in <= 24'b101011111100001111001101;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101001111011101011000100;
#10000;
	data_in <= 24'b101000111011010110111111;
#10000;
	data_in <= 24'b101101111100101111010101;
#10000;
	data_in <= 24'b101101001100101011010100;
#10000;
	data_in <= 24'b101100101100011111010001;
#10000;
	data_in <= 24'b101011101100001111001101;
#10000;
	data_in <= 24'b101010111100000011001010;
#10000;
	data_in <= 24'b101010001011110011000110;
#10000;
	data_in <= 24'b101001011011100011000010;
#10000;
	data_in <= 24'b101000101011010110111111;
#10000;
	data_in <= 24'b110000111100111111010110;
#10000;
	data_in <= 24'b101101101100101111010100;
#10000;
	data_in <= 24'b101100101100100011010010;
#10000;
	data_in <= 24'b101011111100010011001110;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101010011011110011000110;
#10000;
	data_in <= 24'b101001101011100111000011;
#10000;
	data_in <= 24'b101000111011011010111111;
#10000;
	data_in <= 24'b110011101101100011011100;
#10000;
	data_in <= 24'b101111011100110111010101;
#10000;
	data_in <= 24'b101100011100011111010010;
#10000;
	data_in <= 24'b101100001100010011001110;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101010011011110011000110;
#10000;
	data_in <= 24'b101001101011100111000011;
#10000;
	data_in <= 24'b101000101011011010111111;
#10000;
	data_in <= 24'b110100111101110011100001;
#10000;
	data_in <= 24'b110000111101000111011000;
#10000;
	data_in <= 24'b101100011100011111010001;
#10000;
	data_in <= 24'b101011111100001111001101;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101001011011100011000011;
#10000;
	data_in <= 24'b101000111011010110111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100100111010010010101010;
#10000;
	data_in <= 24'b101011101010110010011101;
#10000;
	data_in <= 24'b110100011011111110100000;
#10000;
	data_in <= 24'b110110111100011110101001;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110001100010110100110;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b100000101001011010011111;
#10000;
	data_in <= 24'b110010011011110110100101;
#10000;
	data_in <= 24'b111000001100110010101100;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b100011011010010010110011;
#10000;
	data_in <= 24'b101011111011000110101001;
#10000;
	data_in <= 24'b110111111100101010101010;
#10000;
	data_in <= 24'b110110101100011010101001;
#10000;
	data_in <= 24'b110110011100010110100111;
#10000;
	data_in <= 24'b110110011100010110100111;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b110101111100001110100100;
#10000;
	data_in <= 24'b100101001010100110110110;
#10000;
	data_in <= 24'b100110001010010110101001;
#10000;
	data_in <= 24'b110110011100100010101001;
#10000;
	data_in <= 24'b110110111100100010101001;
#10000;
	data_in <= 24'b110110011100011010100111;
#10000;
	data_in <= 24'b110110011100011010100111;
#10000;
	data_in <= 24'b110101111100010110100101;
#10000;
	data_in <= 24'b110101111100010010100100;
#10000;
	data_in <= 24'b100110011010110110111001;
#10000;
	data_in <= 24'b100011111010000110101011;
#10000;
	data_in <= 24'b110011111100001010101000;
#10000;
	data_in <= 24'b110111011100100110101010;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100001110100100;
#10000;
	data_in <= 24'b100111001010111110111010;
#10000;
	data_in <= 24'b100011001010000110101100;
#10000;
	data_in <= 24'b110001101011110110100111;
#10000;
	data_in <= 24'b110111111100101010101010;
#10000;
	data_in <= 24'b110110001100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100001110100100;
#10000;
	data_in <= 24'b100111001010111110111010;
#10000;
	data_in <= 24'b100010111010000010101100;
#10000;
	data_in <= 24'b110000111011101110101000;
#10000;
	data_in <= 24'b110111111100101010101010;
#10000;
	data_in <= 24'b110110001100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100001110100101;
#10000;
	data_in <= 24'b100111001010111110111010;
#10000;
	data_in <= 24'b100010111010000010101100;
#10000;
	data_in <= 24'b110001001011101110101000;
#10000;
	data_in <= 24'b110111111100101110101010;
#10000;
	data_in <= 24'b110110001100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101011100001010100010;
#10000;
	data_in <= 24'b110100111100000010100000;
#10000;
	data_in <= 24'b110100011011110110011101;
#10000;
	data_in <= 24'b110100001011101110011100;
#10000;
	data_in <= 24'b110011101011101010011001;
#10000;
	data_in <= 24'b110010111011011110010111;
#10000;
	data_in <= 24'b110010011011011010010100;
#10000;
	data_in <= 24'b110001111011001110010010;
#10000;
	data_in <= 24'b110101011100001010100011;
#10000;
	data_in <= 24'b110100111100000010100000;
#10000;
	data_in <= 24'b110100011011110010011101;
#10000;
	data_in <= 24'b110100001011101110011100;
#10000;
	data_in <= 24'b110011101011101010011010;
#10000;
	data_in <= 24'b110010111011011110011000;
#10000;
	data_in <= 24'b110010011011011010010101;
#10000;
	data_in <= 24'b110001101011001110010010;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110101001100000010100000;
#10000;
	data_in <= 24'b110100101011110110011101;
#10000;
	data_in <= 24'b110100011011101110011100;
#10000;
	data_in <= 24'b110011111011101010011011;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110010101011011010010101;
#10000;
	data_in <= 24'b110001111011001110010010;
#10000;
	data_in <= 24'b110101101100001010100010;
#10000;
	data_in <= 24'b110101001100000010100000;
#10000;
	data_in <= 24'b110100101011111010011110;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100001011101110011011;
#10000;
	data_in <= 24'b110011011011100110011000;
#10000;
	data_in <= 24'b110010101011011110010101;
#10000;
	data_in <= 24'b110010001011010010010011;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110101001100000010100001;
#10000;
	data_in <= 24'b110100101011111010011111;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110011111011101110011011;
#10000;
	data_in <= 24'b110011001011100010011000;
#10000;
	data_in <= 24'b110010101011011010010110;
#10000;
	data_in <= 24'b110001111011001110010011;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110101001100000010100001;
#10000;
	data_in <= 24'b110100101011111010011111;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110011111011101110011010;
#10000;
	data_in <= 24'b110011001011100110011000;
#10000;
	data_in <= 24'b110010101011011010010111;
#10000;
	data_in <= 24'b110001111011010010010011;
#10000;
	data_in <= 24'b110101101100001010100011;
#10000;
	data_in <= 24'b110101001100000010100010;
#10000;
	data_in <= 24'b110100101011111010011111;
#10000;
	data_in <= 24'b110100001011110010011101;
#10000;
	data_in <= 24'b110011101011101010011011;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110010101011010110010111;
#10000;
	data_in <= 24'b110001111011001110010100;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110101001100000110100001;
#10000;
	data_in <= 24'b110100101011111110011111;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110011111011101010011100;
#10000;
	data_in <= 24'b110011011011100010011010;
#10000;
	data_in <= 24'b110010101011011010010111;
#10000;
	data_in <= 24'b110001111011010010010100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110000111010110110001110;
#10000;
	data_in <= 24'b110000001010101110001010;
#10000;
	data_in <= 24'b101111011010100010000110;
#10000;
	data_in <= 24'b101110111010011010000100;
#10000;
	data_in <= 24'b101110001010001110000000;
#10000;
	data_in <= 24'b101101001010000001111100;
#10000;
	data_in <= 24'b101100101001110001111010;
#10000;
	data_in <= 24'b110001011010111110010000;
#10000;
	data_in <= 24'b110000111010111010001110;
#10000;
	data_in <= 24'b110000001010101110001010;
#10000;
	data_in <= 24'b101111011010100010000111;
#10000;
	data_in <= 24'b101110111010011010000101;
#10000;
	data_in <= 24'b101110001010001110000001;
#10000;
	data_in <= 24'b101101011001111101111101;
#10000;
	data_in <= 24'b101100101001110001111011;
#10000;
	data_in <= 24'b110001011011000010010000;
#10000;
	data_in <= 24'b110001001010111010001110;
#10000;
	data_in <= 24'b110000011010101110001010;
#10000;
	data_in <= 24'b101111101010100110000111;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101101101001111101111110;
#10000;
	data_in <= 24'b101101001001110001111011;
#10000;
	data_in <= 24'b110001011011001010010000;
#10000;
	data_in <= 24'b110001001010111110001110;
#10000;
	data_in <= 24'b110000011010110010001011;
#10000;
	data_in <= 24'b101111101010100110000111;
#10000;
	data_in <= 24'b101111001010011010000100;
#10000;
	data_in <= 24'b101110011010001110000001;
#10000;
	data_in <= 24'b101101101010000001111110;
#10000;
	data_in <= 24'b101101001001110101111010;
#10000;
	data_in <= 24'b110001011011000110010000;
#10000;
	data_in <= 24'b110001001011000010001110;
#10000;
	data_in <= 24'b110000011010110010001100;
#10000;
	data_in <= 24'b101111101010100110001000;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101101101010000001111110;
#10000;
	data_in <= 24'b101101001001111001111011;
#10000;
	data_in <= 24'b110001011011000110010000;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b101111101010100010001000;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101101101010000001111110;
#10000;
	data_in <= 24'b101101001001111001111011;
#10000;
	data_in <= 24'b110001011011000110010001;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b101111101010100010001001;
#10000;
	data_in <= 24'b101111001010011010000101;
#10000;
	data_in <= 24'b101110011010001110000010;
#10000;
	data_in <= 24'b101101101010000001111111;
#10000;
	data_in <= 24'b101101001001111001111100;
#10000;
	data_in <= 24'b110001011011001010010001;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b101111101010100110001001;
#10000;
	data_in <= 24'b101111001010011010000110;
#10000;
	data_in <= 24'b101110011010010010000010;
#10000;
	data_in <= 24'b101101101010000101111111;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101011111001100101110111;
#10000;
	data_in <= 24'b101010111001010101110010;
#10000;
	data_in <= 24'b101010001001000101101110;
#10000;
	data_in <= 24'b101001001000111001101010;
#10000;
	data_in <= 24'b101000011000101101100110;
#10000;
	data_in <= 24'b100111011000011101100011;
#10000;
	data_in <= 24'b100110101000001101011110;
#10000;
	data_in <= 24'b100101010111110101011010;
#10000;
	data_in <= 24'b101011101001100001110111;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101001111001000101101111;
#10000;
	data_in <= 24'b101001001000111001101011;
#10000;
	data_in <= 24'b101000011000101001100111;
#10000;
	data_in <= 24'b100111011000011101100011;
#10000;
	data_in <= 24'b100110101000001001011111;
#10000;
	data_in <= 24'b100101100111110101011011;
#10000;
	data_in <= 24'b101100001001100101110110;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101010001001001001101111;
#10000;
	data_in <= 24'b101001011000111001101011;
#10000;
	data_in <= 24'b101000011000101101101000;
#10000;
	data_in <= 24'b100111101000011101100100;
#10000;
	data_in <= 24'b100110101000001001100000;
#10000;
	data_in <= 24'b100101100111111001011100;
#10000;
	data_in <= 24'b101100001001101001110110;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101010001001001001101111;
#10000;
	data_in <= 24'b101001011000111101101011;
#10000;
	data_in <= 24'b101000101000110001100111;
#10000;
	data_in <= 24'b100111101000100001100011;
#10000;
	data_in <= 24'b100110111000010001011111;
#10000;
	data_in <= 24'b100101101000000001011011;
#10000;
	data_in <= 24'b101100001001100101110111;
#10000;
	data_in <= 24'b101010111001010101110100;
#10000;
	data_in <= 24'b101010001001001001110000;
#10000;
	data_in <= 24'b101001011000111101101100;
#10000;
	data_in <= 24'b101000011000101101101000;
#10000;
	data_in <= 24'b100111101000011101100100;
#10000;
	data_in <= 24'b100110111000001101100000;
#10000;
	data_in <= 24'b100101100111111101011011;
#10000;
	data_in <= 24'b101011111001100101111000;
#10000;
	data_in <= 24'b101010111001010101110011;
#10000;
	data_in <= 24'b101010001001001001101111;
#10000;
	data_in <= 24'b101001011000111101101101;
#10000;
	data_in <= 24'b101000011000101101101001;
#10000;
	data_in <= 24'b100111101000011101100100;
#10000;
	data_in <= 24'b100110111000010001100000;
#10000;
	data_in <= 24'b100101100111111101011011;
#10000;
	data_in <= 24'b101011111001100101111000;
#10000;
	data_in <= 24'b101010111001010101110100;
#10000;
	data_in <= 24'b101010001001001001110001;
#10000;
	data_in <= 24'b101001011000111101101101;
#10000;
	data_in <= 24'b101000011000101101101001;
#10000;
	data_in <= 24'b100111101000011101100101;
#10000;
	data_in <= 24'b100110111000001101100001;
#10000;
	data_in <= 24'b100101100111111101011100;
#10000;
	data_in <= 24'b101100001001101001111001;
#10000;
	data_in <= 24'b101010111001011001110100;
#10000;
	data_in <= 24'b101010001001001001110010;
#10000;
	data_in <= 24'b101001011001000001101101;
#10000;
	data_in <= 24'b101000011000101101101001;
#10000;
	data_in <= 24'b100111101000011101100110;
#10000;
	data_in <= 24'b100110111000010001100010;
#10000;
	data_in <= 24'b100101101000000001011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100101101000000101011110;
#10000;
	data_in <= 24'b100110111000010101100010;
#10000;
	data_in <= 24'b100111101000100001100110;
#10000;
	data_in <= 24'b101000101000101101101010;
#10000;
	data_in <= 24'b101001011001000001101101;
#10000;
	data_in <= 24'b101010001001001101110001;
#10000;
	data_in <= 24'b101011001001011101110100;
#10000;
	data_in <= 24'b101011111001101101111000;
#10000;
	data_in <= 24'b100101101000000101011111;
#10000;
	data_in <= 24'b100110111000010101100011;
#10000;
	data_in <= 24'b100111101000100001100111;
#10000;
	data_in <= 24'b101000101000101101101011;
#10000;
	data_in <= 24'b101001011000111101101110;
#10000;
	data_in <= 24'b101010001001010001110010;
#10000;
	data_in <= 24'b101011001001011101110110;
#10000;
	data_in <= 24'b101100001001101001111001;
#10000;
	data_in <= 24'b100101111000000001011110;
#10000;
	data_in <= 24'b100110111000010001100010;
#10000;
	data_in <= 24'b100111101000100001100110;
#10000;
	data_in <= 24'b101000011000101101101010;
#10000;
	data_in <= 24'b101001011000111101101110;
#10000;
	data_in <= 24'b101010011001010001110001;
#10000;
	data_in <= 24'b101011001001011101110110;
#10000;
	data_in <= 24'b101011111001101001111010;
#10000;
	data_in <= 24'b100101101000000001011110;
#10000;
	data_in <= 24'b100110111000010001100010;
#10000;
	data_in <= 24'b100111111000100001100110;
#10000;
	data_in <= 24'b101000111000110101101010;
#10000;
	data_in <= 24'b101001101001000001101110;
#10000;
	data_in <= 24'b101010011001010001110010;
#10000;
	data_in <= 24'b101011001001011101110110;
#10000;
	data_in <= 24'b101100001001101101111010;
#10000;
	data_in <= 24'b100101111000000001011110;
#10000;
	data_in <= 24'b100111001000010101100011;
#10000;
	data_in <= 24'b101000001000101001100111;
#10000;
	data_in <= 24'b101001001000111001101010;
#10000;
	data_in <= 24'b101001111001000101101110;
#10000;
	data_in <= 24'b101010101001010001110011;
#10000;
	data_in <= 24'b101011011001011101110111;
#10000;
	data_in <= 24'b101100011001110001111011;
#10000;
	data_in <= 24'b100110001000000001011110;
#10000;
	data_in <= 24'b100111001000010001100011;
#10000;
	data_in <= 24'b101000001000100101100111;
#10000;
	data_in <= 24'b101001001000111001101011;
#10000;
	data_in <= 24'b101001111001000101101111;
#10000;
	data_in <= 24'b101010101001010001110011;
#10000;
	data_in <= 24'b101011011001011101110110;
#10000;
	data_in <= 24'b101100001001101101111001;
#10000;
	data_in <= 24'b100101111000000101011111;
#10000;
	data_in <= 24'b100110111000010101100011;
#10000;
	data_in <= 24'b101000001000100101101000;
#10000;
	data_in <= 24'b101001001000111001101100;
#10000;
	data_in <= 24'b101001111001000101101111;
#10000;
	data_in <= 24'b101010101001010001110010;
#10000;
	data_in <= 24'b101011011001011101110110;
#10000;
	data_in <= 24'b101100011001101001111010;
#10000;
	data_in <= 24'b100110001000001001100001;
#10000;
	data_in <= 24'b100111001000010101100101;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b101001001000111001101101;
#10000;
	data_in <= 24'b101001111001000101110000;
#10000;
	data_in <= 24'b101010101001010001110011;
#10000;
	data_in <= 24'b101011011001011101110111;
#10000;
	data_in <= 24'b101100011001101001111100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b101101101010000101111111;
#10000;
	data_in <= 24'b101110011010010010000011;
#10000;
	data_in <= 24'b101111001010011110000111;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110001011011001010010010;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b101101101010000110000000;
#10000;
	data_in <= 24'b101110011010010010000100;
#10000;
	data_in <= 24'b101111001010011110000111;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b110000011010110110001101;
#10000;
	data_in <= 24'b110001001011000010010000;
#10000;
	data_in <= 24'b110001011011000110010010;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b101101011010000010000000;
#10000;
	data_in <= 24'b101110011010010010000100;
#10000;
	data_in <= 24'b101111001010011110000111;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b110000011010110110001101;
#10000;
	data_in <= 24'b110001001011000010010000;
#10000;
	data_in <= 24'b110001011011000110010010;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b101101101010000110000000;
#10000;
	data_in <= 24'b101110011010010010000100;
#10000;
	data_in <= 24'b101111001010100010000111;
#10000;
	data_in <= 24'b101111101010101110001001;
#10000;
	data_in <= 24'b110000101010110110001101;
#10000;
	data_in <= 24'b110001001011000010010000;
#10000;
	data_in <= 24'b110001111011001010010011;
#10000;
	data_in <= 24'b101101001001111101111110;
#10000;
	data_in <= 24'b101101101010000110000001;
#10000;
	data_in <= 24'b101110011010010110000100;
#10000;
	data_in <= 24'b101111001010100010001000;
#10000;
	data_in <= 24'b101111101010101110001010;
#10000;
	data_in <= 24'b110000011010111010001101;
#10000;
	data_in <= 24'b110001011011000110010001;
#10000;
	data_in <= 24'b110010001011001110010011;
#10000;
	data_in <= 24'b101101001001111101111110;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101110011010010110000100;
#10000;
	data_in <= 24'b101111001010100010000111;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b110000011010111010001110;
#10000;
	data_in <= 24'b110001001011000110010001;
#10000;
	data_in <= 24'b110001111011001010010010;
#10000;
	data_in <= 24'b101101001001111001111110;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101110011010010110000100;
#10000;
	data_in <= 24'b101111001010100010000111;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b110000011010110110001110;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110001111011001010010011;
#10000;
	data_in <= 24'b101101001001111001111111;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101110011010010110000101;
#10000;
	data_in <= 24'b101111001010100010001000;
#10000;
	data_in <= 24'b101111101010101010001011;
#10000;
	data_in <= 24'b110000011010110110001111;
#10000;
	data_in <= 24'b110001011011000010010010;
#10000;
	data_in <= 24'b110001101011001010010011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110010001011010010010101;
#10000;
	data_in <= 24'b110010111011011110010111;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110011111011101010011011;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110101001100000110100001;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110010001011010010010101;
#10000;
	data_in <= 24'b110010111011011110011000;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110011111011101010011011;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110100011011111010100000;
#10000;
	data_in <= 24'b110100111100000010100010;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110010001011010010010101;
#10000;
	data_in <= 24'b110010111011011010010111;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110011111011101110011100;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100111100000010100010;
#10000;
	data_in <= 24'b110101011100001010100100;
#10000;
	data_in <= 24'b110010011011010010010101;
#10000;
	data_in <= 24'b110010111011011010010111;
#10000;
	data_in <= 24'b110011011011100110011001;
#10000;
	data_in <= 24'b110011111011101110011100;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100111100000010100001;
#10000;
	data_in <= 24'b110101011100001010100100;
#10000;
	data_in <= 24'b110010101011010110010110;
#10000;
	data_in <= 24'b110011001011011110011000;
#10000;
	data_in <= 24'b110011101011100110011010;
#10000;
	data_in <= 24'b110100001011110010011100;
#10000;
	data_in <= 24'b110100011011111010011110;
#10000;
	data_in <= 24'b110100101011111110100000;
#10000;
	data_in <= 24'b110101001100000110100010;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110010101011010010010101;
#10000;
	data_in <= 24'b110010111011011110011000;
#10000;
	data_in <= 24'b110011011011100110011010;
#10000;
	data_in <= 24'b110100001011110010011101;
#10000;
	data_in <= 24'b110100011011111010011110;
#10000;
	data_in <= 24'b110100101011111110011111;
#10000;
	data_in <= 24'b110101001100000110100010;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b110010011011010010010101;
#10000;
	data_in <= 24'b110011001011011110011000;
#10000;
	data_in <= 24'b110011011011100110011011;
#10000;
	data_in <= 24'b110100001011101110011101;
#10000;
	data_in <= 24'b110100011011110110011110;
#10000;
	data_in <= 24'b110100101011111110011111;
#10000;
	data_in <= 24'b110101001100000110100010;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b110010011011010110010110;
#10000;
	data_in <= 24'b110011001011011110011001;
#10000;
	data_in <= 24'b110011011011100110011100;
#10000;
	data_in <= 24'b110100001011110010011110;
#10000;
	data_in <= 24'b110100011011110110011111;
#10000;
	data_in <= 24'b110100101011111010100000;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110111100100110101010;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101001;
#10000;
	data_in <= 24'b110110111100100110101011;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b110110001100010010100110;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011110101000;
#10000;
	data_in <= 24'b110110101100100110101010;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110101101100001110100110;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011110101000;
#10000;
	data_in <= 24'b110110111100100110101010;
#10000;
	data_in <= 24'b110111001100101010101011;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100010010101000;
#10000;
	data_in <= 24'b110110011100011010101001;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110110111100100110101011;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110110011100011010101001;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110110011100011110101000;
#10000;
	data_in <= 24'b110110101100011110101010;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110110101100011110101010;
#10000;
	data_in <= 24'b110111001100100010101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110111101100110010101110;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b110111101100110110101111;
#10000;
	data_in <= 24'b111000001100111010101110;
#10000;
	data_in <= 24'b101000011010101010101000;
#10000;
	data_in <= 24'b100011011010010010110010;
#10000;
	data_in <= 24'b101000001011001110111100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b110111101100110010110000;
#10000;
	data_in <= 24'b110111011100110010110000;
#10000;
	data_in <= 24'b111001001101000010110001;
#10000;
	data_in <= 24'b101011101011000110101000;
#10000;
	data_in <= 24'b100010101010000010101110;
#10000;
	data_in <= 24'b100111111011000110111011;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b110111001100101110101111;
#10000;
	data_in <= 24'b111001001101000010110001;
#10000;
	data_in <= 24'b110001011011111010101010;
#10000;
	data_in <= 24'b100010011001111010101001;
#10000;
	data_in <= 24'b100110011010110010111000;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110111101100101110101111;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111101100110110101111;
#10000;
	data_in <= 24'b100110001010010010100101;
#10000;
	data_in <= 24'b100011101010010010110001;
#10000;
	data_in <= 24'b110111101100101110101110;
#10000;
	data_in <= 24'b110111111100110010110000;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111101100110010110000;
#10000;
	data_in <= 24'b111001001101000010110001;
#10000;
	data_in <= 24'b110000111011110010101010;
#10000;
	data_in <= 24'b100001101001110010100111;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b111001001101000010110001;
#10000;
	data_in <= 24'b101010111010111110100111;
#10000;
	data_in <= 24'b110111011100101010101110;
#10000;
	data_in <= 24'b110111101100110010101111;
#10000;
	data_in <= 24'b110111101100110110101111;
#10000;
	data_in <= 24'b110111101100110110101111;
#10000;
	data_in <= 24'b110111101100110110101111;
#10000;
	data_in <= 24'b110111101100110110110000;
#10000;
	data_in <= 24'b110111111100110110110000;
#10000;
	data_in <= 24'b111000011100111010110001;
#10000;
	data_in <= 24'b110111011100101010101110;
#10000;
	data_in <= 24'b110111101100101110110000;
#10000;
	data_in <= 24'b110111101100110010110000;
#10000;
	data_in <= 24'b110111101100110010110000;
#10000;
	data_in <= 24'b110111011100110010110000;
#10000;
	data_in <= 24'b110111101100110110110000;
#10000;
	data_in <= 24'b111000101101000010110000;
#10000;
	data_in <= 24'b110111111100110110110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000111011011011000000;
#10000;
	data_in <= 24'b101001101011100111000100;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101011111100010011001110;
#10000;
	data_in <= 24'b101101001100100011010010;
#10000;
	data_in <= 24'b110010111101011111011100;
#10000;
	data_in <= 24'b110101001101111011100011;
#10000;
	data_in <= 24'b101000101011010110111111;
#10000;
	data_in <= 24'b101001011011100111000011;
#10000;
	data_in <= 24'b101010001011110011000110;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101011011100001011001100;
#10000;
	data_in <= 24'b101100111100011111010001;
#10000;
	data_in <= 24'b110010111101011111011100;
#10000;
	data_in <= 24'b110101011101111111100100;
#10000;
	data_in <= 24'b101000011011010010111110;
#10000;
	data_in <= 24'b101001001011011111000010;
#10000;
	data_in <= 24'b101001111011101011000101;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101100011100010111001111;
#10000;
	data_in <= 24'b110010101101011011011100;
#10000;
	data_in <= 24'b110101011101111011100011;
#10000;
	data_in <= 24'b101000001011001010111100;
#10000;
	data_in <= 24'b101000111011010111000000;
#10000;
	data_in <= 24'b101001011011100111000011;
#10000;
	data_in <= 24'b101010001011110011000110;
#10000;
	data_in <= 24'b101010111011111111001001;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b110000111101000011011000;
#10000;
	data_in <= 24'b110101011101111011100010;
#10000;
	data_in <= 24'b100110001010110010110110;
#10000;
	data_in <= 24'b101000011011010010111110;
#10000;
	data_in <= 24'b101000111011011011000001;
#10000;
	data_in <= 24'b101001101011101011000100;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101101001100011011001111;
#10000;
	data_in <= 24'b110100001101101011011111;
#10000;
	data_in <= 24'b100000111001110010101010;
#10000;
	data_in <= 24'b100110101010110110111000;
#10000;
	data_in <= 24'b101000011011010010111110;
#10000;
	data_in <= 24'b101001001011011111000001;
#10000;
	data_in <= 24'b101001111011101011000100;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101010011011111011001000;
#10000;
	data_in <= 24'b101111001100110011010100;
#10000;
	data_in <= 24'b101010111010111010100111;
#10000;
	data_in <= 24'b100011001010000010101010;
#10000;
	data_in <= 24'b100110011010110110110111;
#10000;
	data_in <= 24'b101000001011010010111110;
#10000;
	data_in <= 24'b101001001011011111000001;
#10000;
	data_in <= 24'b101001101011101011000100;
#10000;
	data_in <= 24'b101010001011110011000110;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b110001011011111110101101;
#10000;
	data_in <= 24'b100010101001110010100010;
#10000;
	data_in <= 24'b100001101001101110100110;
#10000;
	data_in <= 24'b100101011010100010110010;
#10000;
	data_in <= 24'b100111011011000010111011;
#10000;
	data_in <= 24'b101000101011010110111111;
#10000;
	data_in <= 24'b101001011011100011000010;
#10000;
	data_in <= 24'b101001111011101011000101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101111110001011100110;
#10000;
	data_in <= 24'b110110101110010111101010;
#10000;
	data_in <= 24'b110111101110100111101101;
#10000;
	data_in <= 24'b111000001110101111101111;
#10000;
	data_in <= 24'b110111111110101111101111;
#10000;
	data_in <= 24'b110111101110100111101110;
#10000;
	data_in <= 24'b110110101110011011101010;
#10000;
	data_in <= 24'b110101111110000111100111;
#10000;
	data_in <= 24'b110101111110001011100110;
#10000;
	data_in <= 24'b110110101110011011101011;
#10000;
	data_in <= 24'b110111111110101011101111;
#10000;
	data_in <= 24'b111000011110110111110001;
#10000;
	data_in <= 24'b111000011110110011110001;
#10000;
	data_in <= 24'b110111101110100111101111;
#10000;
	data_in <= 24'b110110111110011011101011;
#10000;
	data_in <= 24'b110101111110001011100111;
#10000;
	data_in <= 24'b110101111110000111100110;
#10000;
	data_in <= 24'b110110101110010111101010;
#10000;
	data_in <= 24'b110111011110100111101101;
#10000;
	data_in <= 24'b110111111110101111101111;
#10000;
	data_in <= 24'b110111111110101111110000;
#10000;
	data_in <= 24'b110111101110100111101110;
#10000;
	data_in <= 24'b110110101110010111101010;
#10000;
	data_in <= 24'b110101111110001011100111;
#10000;
	data_in <= 24'b110101011110000011100101;
#10000;
	data_in <= 24'b110110011110001111101000;
#10000;
	data_in <= 24'b110110111110011011101011;
#10000;
	data_in <= 24'b110111001110011111101100;
#10000;
	data_in <= 24'b110111001110100011101100;
#10000;
	data_in <= 24'b110110111110011011101011;
#10000;
	data_in <= 24'b110110001110001111101000;
#10000;
	data_in <= 24'b110101101110000011100101;
#10000;
	data_in <= 24'b110101001101111011100011;
#10000;
	data_in <= 24'b110101011110000011100101;
#10000;
	data_in <= 24'b110110001110001011100111;
#10000;
	data_in <= 24'b110110011110001111101001;
#10000;
	data_in <= 24'b110110011110010011101000;
#10000;
	data_in <= 24'b110101111110001011100111;
#10000;
	data_in <= 24'b110101011110000011100101;
#10000;
	data_in <= 24'b110101101101111111100100;
#10000;
	data_in <= 24'b110100111101110011100001;
#10000;
	data_in <= 24'b110101011101111111100011;
#10000;
	data_in <= 24'b110101011101111111100100;
#10000;
	data_in <= 24'b110101011101111111100100;
#10000;
	data_in <= 24'b110101011101111111100100;
#10000;
	data_in <= 24'b110101011101111111100100;
#10000;
	data_in <= 24'b110101101101111111100011;
#10000;
	data_in <= 24'b110011101101100111011110;
#10000;
	data_in <= 24'b101110011100100111010001;
#10000;
	data_in <= 24'b110011001101011111011101;
#10000;
	data_in <= 24'b110100111101110011100001;
#10000;
	data_in <= 24'b110101011101111011100011;
#10000;
	data_in <= 24'b110101011101111011100011;
#10000;
	data_in <= 24'b110100101101101111100001;
#10000;
	data_in <= 24'b110010001101010011011010;
#10000;
	data_in <= 24'b101100011100001111001100;
#10000;
	data_in <= 24'b101001101011101011000101;
#10000;
	data_in <= 24'b101010111011111111001001;
#10000;
	data_in <= 24'b101101011100011011001111;
#10000;
	data_in <= 24'b101111011100110011010011;
#10000;
	data_in <= 24'b101111001100101111010011;
#10000;
	data_in <= 24'b101100111100010011001101;
#10000;
	data_in <= 24'b101010001011110011000110;
#10000;
	data_in <= 24'b101001101011101011000100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101001101111011100011;
#10000;
	data_in <= 24'b110001111101001111011010;
#10000;
	data_in <= 24'b101100011100011011010000;
#10000;
	data_in <= 24'b101011101100001111001101;
#10000;
	data_in <= 24'b101010111011111111001001;
#10000;
	data_in <= 24'b101010001011101111000110;
#10000;
	data_in <= 24'b101001011011100011000010;
#10000;
	data_in <= 24'b101000101011010110111110;
#10000;
	data_in <= 24'b110101011101111111100011;
#10000;
	data_in <= 24'b110001111101001111011001;
#10000;
	data_in <= 24'b101011111100010011001110;
#10000;
	data_in <= 24'b101011011100001011001100;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101001111011101011000101;
#10000;
	data_in <= 24'b101001001011011111000001;
#10000;
	data_in <= 24'b101000011011010010111110;
#10000;
	data_in <= 24'b110101011101111011100011;
#10000;
	data_in <= 24'b110000001101000011010111;
#10000;
	data_in <= 24'b101011001100001011001101;
#10000;
	data_in <= 24'b101011001100000011001010;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101001101011100111000011;
#10000;
	data_in <= 24'b101000111011011011000000;
#10000;
	data_in <= 24'b101000001011001010111100;
#10000;
	data_in <= 24'b110100101101110011100001;
#10000;
	data_in <= 24'b101101111100100111010010;
#10000;
	data_in <= 24'b101010111100000011001010;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101001111011101111000101;
#10000;
	data_in <= 24'b101001001011100011000010;
#10000;
	data_in <= 24'b101000101011010010111110;
#10000;
	data_in <= 24'b100110101010110110111001;
#10000;
	data_in <= 24'b110010001101010011011010;
#10000;
	data_in <= 24'b101011001100000111001011;
#10000;
	data_in <= 24'b101010101011111011001000;
#10000;
	data_in <= 24'b101010001011101111000101;
#10000;
	data_in <= 24'b101001011011100111000011;
#10000;
	data_in <= 24'b101000111011011011000000;
#10000;
	data_in <= 24'b100111101011000110111011;
#10000;
	data_in <= 24'b100010001010000110101110;
#10000;
	data_in <= 24'b101100101100010011001110;
#10000;
	data_in <= 24'b101010011011110111000111;
#10000;
	data_in <= 24'b101010001011101111000110;
#10000;
	data_in <= 24'b101001101011100111000100;
#10000;
	data_in <= 24'b101000111011011011000000;
#10000;
	data_in <= 24'b100111111011001010111100;
#10000;
	data_in <= 24'b100100101010011110110010;
#10000;
	data_in <= 24'b100101101010001110100110;
#10000;
	data_in <= 24'b101010001011110011000110;
#10000;
	data_in <= 24'b101010001011110011000110;
#10000;
	data_in <= 24'b101001101011100111000011;
#10000;
	data_in <= 24'b101000101011011011000000;
#10000;
	data_in <= 24'b100111011011000110111011;
#10000;
	data_in <= 24'b100100111010011110110001;
#10000;
	data_in <= 24'b011111111001011010100001;
#10000;
	data_in <= 24'b101010111010110010100010;
#10000;
	data_in <= 24'b101001101011100111000100;
#10000;
	data_in <= 24'b101000111011011111000001;
#10000;
	data_in <= 24'b100111111011001110111101;
#10000;
	data_in <= 24'b100110001010110010110110;
#10000;
	data_in <= 24'b100011101010001010101100;
#10000;
	data_in <= 24'b100000111001100110100010;
#10000;
	data_in <= 24'b011110011001010010100000;
#10000;
	data_in <= 24'b011100001000111010011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100110101010110110111001;
#10000;
	data_in <= 24'b100011001001111110101010;
#10000;
	data_in <= 24'b110010101011111110101000;
#10000;
	data_in <= 24'b110111101100101010101010;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b100101011010101010110110;
#10000;
	data_in <= 24'b100100011010000110100111;
#10000;
	data_in <= 24'b110101101100010110101010;
#10000;
	data_in <= 24'b110111001100100110101011;
#10000;
	data_in <= 24'b110110011100011010101001;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101111100010010100101;
#10000;
	data_in <= 24'b100011001010001110110000;
#10000;
	data_in <= 24'b101000111010101010100110;
#10000;
	data_in <= 24'b110111111100101110101100;
#10000;
	data_in <= 24'b110110101100100110101010;
#10000;
	data_in <= 24'b110110011100011110101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110001100010010100110;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b100001111001110110101000;
#10000;
	data_in <= 24'b110001001011101110101000;
#10000;
	data_in <= 24'b111000011100110010101100;
#10000;
	data_in <= 24'b110110101100100110101010;
#10000;
	data_in <= 24'b110110011100011110101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101101100001110100110;
#10000;
	data_in <= 24'b101000001010100010100101;
#10000;
	data_in <= 24'b110111101100101110101100;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110110101100100010101011;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110101111100010010101000;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100011010101100;
#10000;
	data_in <= 24'b111000101100110110101110;
#10000;
	data_in <= 24'b110110111100100110101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110110011100011010101001;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110110001100011110101100;
#10000;
	data_in <= 24'b110110101100100010101100;
#10000;
	data_in <= 24'b110111111100101010101100;
#10000;
	data_in <= 24'b111000001100101110101100;
#10000;
	data_in <= 24'b110111101100100110101010;
#10000;
	data_in <= 24'b110111011100100110101001;
#10000;
	data_in <= 24'b110111011100100010101000;
#10000;
	data_in <= 24'b110111111100100010101000;
#10000;
	data_in <= 24'b011100101000110110011000;
#10000;
	data_in <= 24'b011111001001001010011000;
#10000;
	data_in <= 24'b100001001001011110011010;
#10000;
	data_in <= 24'b100001101001100010011011;
#10000;
	data_in <= 24'b100001101001011110011001;
#10000;
	data_in <= 24'b100001111001011110011000;
#10000;
	data_in <= 24'b100011011001101010011000;
#10000;
	data_in <= 24'b100110001001111110011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110101001100000110100001;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110011111011101010011011;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110010111011011110010111;
#10000;
	data_in <= 24'b110010001011010010010101;
#10000;
	data_in <= 24'b110101101100001110100011;
#10000;
	data_in <= 24'b110100111100000010100010;
#10000;
	data_in <= 24'b110100011011111010100000;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110011111011101010011011;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110010111011011110011000;
#10000;
	data_in <= 24'b110010001011010010010101;
#10000;
	data_in <= 24'b110101011100001010100100;
#10000;
	data_in <= 24'b110100111100000010100010;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110011111011101110011100;
#10000;
	data_in <= 24'b110011001011100010011001;
#10000;
	data_in <= 24'b110010111011011010010111;
#10000;
	data_in <= 24'b110010001011010010010101;
#10000;
	data_in <= 24'b110101011100001010100100;
#10000;
	data_in <= 24'b110100111100000010100001;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100001011110110011110;
#10000;
	data_in <= 24'b110011111011101110011100;
#10000;
	data_in <= 24'b110011011011100110011001;
#10000;
	data_in <= 24'b110010111011011010010111;
#10000;
	data_in <= 24'b110010011011010010010101;
#10000;
	data_in <= 24'b110101101100001110100100;
#10000;
	data_in <= 24'b110101001100000110100010;
#10000;
	data_in <= 24'b110100101011111110100000;
#10000;
	data_in <= 24'b110100011011111010011110;
#10000;
	data_in <= 24'b110100001011110010011100;
#10000;
	data_in <= 24'b110011101011100110011010;
#10000;
	data_in <= 24'b110011001011011110011000;
#10000;
	data_in <= 24'b110010101011010110010110;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110100101100000010100010;
#10000;
	data_in <= 24'b110100101011111110011111;
#10000;
	data_in <= 24'b110100011011111010011110;
#10000;
	data_in <= 24'b110100001011110010011101;
#10000;
	data_in <= 24'b110011011011100110011010;
#10000;
	data_in <= 24'b110011001011011110011000;
#10000;
	data_in <= 24'b110010101011010010010101;
#10000;
	data_in <= 24'b110111111100100010100111;
#10000;
	data_in <= 24'b110110101100010110100011;
#10000;
	data_in <= 24'b110100111011111110011111;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110011111011101110011101;
#10000;
	data_in <= 24'b110011011011101010011011;
#10000;
	data_in <= 24'b110011001011011110011000;
#10000;
	data_in <= 24'b110010011011010010010101;
#10000;
	data_in <= 24'b101010001010100010011011;
#10000;
	data_in <= 24'b101111101011010010011110;
#10000;
	data_in <= 24'b110101001011111110100000;
#10000;
	data_in <= 24'b110110011100000110100000;
#10000;
	data_in <= 24'b110100001011110010011110;
#10000;
	data_in <= 24'b110011011011100110011011;
#10000;
	data_in <= 24'b110011001011011110011001;
#10000;
	data_in <= 24'b110010011011010110010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001011011001010010010;
#10000;
	data_in <= 24'b110001001011000010001111;
#10000;
	data_in <= 24'b110000011010110110001100;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b101111001010011110000111;
#10000;
	data_in <= 24'b101110011010010010000011;
#10000;
	data_in <= 24'b101101101010000101111111;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b110001011011000110010010;
#10000;
	data_in <= 24'b110001001011000010010000;
#10000;
	data_in <= 24'b110000011010110110001101;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b101111001010011110000111;
#10000;
	data_in <= 24'b101110011010010010000100;
#10000;
	data_in <= 24'b101101101010000110000000;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b110001011011000110010010;
#10000;
	data_in <= 24'b110001001011000010010000;
#10000;
	data_in <= 24'b110000011010110110001101;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b101111001010011110000111;
#10000;
	data_in <= 24'b101110011010010010000100;
#10000;
	data_in <= 24'b101101011010000010000000;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b110001111011001010010011;
#10000;
	data_in <= 24'b110001001011000010010000;
#10000;
	data_in <= 24'b110000101010110110001101;
#10000;
	data_in <= 24'b101111101010101110001001;
#10000;
	data_in <= 24'b101111001010100010000111;
#10000;
	data_in <= 24'b101110011010010010000100;
#10000;
	data_in <= 24'b101101101010000110000000;
#10000;
	data_in <= 24'b101100111001111001111101;
#10000;
	data_in <= 24'b110010001011001110010011;
#10000;
	data_in <= 24'b110001011011000110010001;
#10000;
	data_in <= 24'b110000011010111010001101;
#10000;
	data_in <= 24'b101111101010101110001010;
#10000;
	data_in <= 24'b101111001010100010001000;
#10000;
	data_in <= 24'b101110011010010110000100;
#10000;
	data_in <= 24'b101101101010000110000001;
#10000;
	data_in <= 24'b101101001001111101111110;
#10000;
	data_in <= 24'b110001111011001010010010;
#10000;
	data_in <= 24'b110001001011000110010001;
#10000;
	data_in <= 24'b110000011010111010001110;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b101111001010100010000111;
#10000;
	data_in <= 24'b101110011010010110000100;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101101001001111101111110;
#10000;
	data_in <= 24'b110001111011001010010011;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110000011010110110001110;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b101111001010100010000111;
#10000;
	data_in <= 24'b101110011010010110000100;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101101001001111001111110;
#10000;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b110001011011000010010010;
#10000;
	data_in <= 24'b110000011010110110001111;
#10000;
	data_in <= 24'b101111101010101010001011;
#10000;
	data_in <= 24'b101111001010100010001000;
#10000;
	data_in <= 24'b101110011010010110000101;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101101001001111001111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101011111001101101111000;
#10000;
	data_in <= 24'b101011001001011101110100;
#10000;
	data_in <= 24'b101010001001001101110001;
#10000;
	data_in <= 24'b101001011001000001101101;
#10000;
	data_in <= 24'b101000101000101101101010;
#10000;
	data_in <= 24'b100111101000100001100110;
#10000;
	data_in <= 24'b100110111000010101100010;
#10000;
	data_in <= 24'b100101101000000101011110;
#10000;
	data_in <= 24'b101100001001101001111001;
#10000;
	data_in <= 24'b101011001001011101110110;
#10000;
	data_in <= 24'b101010001001010001110010;
#10000;
	data_in <= 24'b101001011000111101101110;
#10000;
	data_in <= 24'b101000101000101101101011;
#10000;
	data_in <= 24'b100111101000100001100111;
#10000;
	data_in <= 24'b100110111000010101100011;
#10000;
	data_in <= 24'b100101101000000101011111;
#10000;
	data_in <= 24'b101011111001101001111010;
#10000;
	data_in <= 24'b101011001001011101110110;
#10000;
	data_in <= 24'b101010011001010001110001;
#10000;
	data_in <= 24'b101001011000111101101110;
#10000;
	data_in <= 24'b101000011000101101101010;
#10000;
	data_in <= 24'b100111101000100001100110;
#10000;
	data_in <= 24'b100110111000010001100010;
#10000;
	data_in <= 24'b100101111000000001011110;
#10000;
	data_in <= 24'b101100001001101101111010;
#10000;
	data_in <= 24'b101011001001011101110110;
#10000;
	data_in <= 24'b101010011001010001110010;
#10000;
	data_in <= 24'b101001101001000001101110;
#10000;
	data_in <= 24'b101000111000110101101010;
#10000;
	data_in <= 24'b100111111000100001100110;
#10000;
	data_in <= 24'b100110111000010001100010;
#10000;
	data_in <= 24'b100101101000000001011110;
#10000;
	data_in <= 24'b101100011001110001111011;
#10000;
	data_in <= 24'b101011011001011101110111;
#10000;
	data_in <= 24'b101010101001010001110011;
#10000;
	data_in <= 24'b101001111001000101101110;
#10000;
	data_in <= 24'b101001001000111001101010;
#10000;
	data_in <= 24'b101000001000101001100111;
#10000;
	data_in <= 24'b100111001000010101100011;
#10000;
	data_in <= 24'b100101111000000001011110;
#10000;
	data_in <= 24'b101100001001101101111001;
#10000;
	data_in <= 24'b101011011001011101110110;
#10000;
	data_in <= 24'b101010101001010001110011;
#10000;
	data_in <= 24'b101001111001000101101111;
#10000;
	data_in <= 24'b101001001000111001101011;
#10000;
	data_in <= 24'b101000001000100101100111;
#10000;
	data_in <= 24'b100111001000010001100011;
#10000;
	data_in <= 24'b100110001000000001011110;
#10000;
	data_in <= 24'b101100011001101001111010;
#10000;
	data_in <= 24'b101011011001011101110110;
#10000;
	data_in <= 24'b101010101001010001110010;
#10000;
	data_in <= 24'b101001111001000101101111;
#10000;
	data_in <= 24'b101001001000111001101100;
#10000;
	data_in <= 24'b101000001000100101101000;
#10000;
	data_in <= 24'b100110111000010101100011;
#10000;
	data_in <= 24'b100101111000000101011111;
#10000;
	data_in <= 24'b101100011001101001111100;
#10000;
	data_in <= 24'b101011011001011101110111;
#10000;
	data_in <= 24'b101010101001010001110011;
#10000;
	data_in <= 24'b101001111001000101110000;
#10000;
	data_in <= 24'b101001001000111001101101;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b100111001000010101100101;
#10000;
	data_in <= 24'b100110001000001001100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b100110111000011001100100;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b101000111000110101101100;
#10000;
	data_in <= 24'b101001111001000101110000;
#10000;
	data_in <= 24'b101010101001010101110011;
#10000;
	data_in <= 24'b101011011001100001110111;
#10000;
	data_in <= 24'b101100001001101101111100;
#10000;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b100110111000011001100100;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b101000101000110101101011;
#10000;
	data_in <= 24'b101001111001000101110000;
#10000;
	data_in <= 24'b101010101001010101110100;
#10000;
	data_in <= 24'b101011011001100101111000;
#10000;
	data_in <= 24'b101100001001110001111011;
#10000;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b100110101000010101100100;
#10000;
	data_in <= 24'b100111111000101001101001;
#10000;
	data_in <= 24'b101000101000110101101101;
#10000;
	data_in <= 24'b101001101001000001110001;
#10000;
	data_in <= 24'b101010101001010001110101;
#10000;
	data_in <= 24'b101011011001100101111000;
#10000;
	data_in <= 24'b101100001001110001111011;
#10000;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b100110101000010101100011;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b101000011000110001101101;
#10000;
	data_in <= 24'b101001101001000101110001;
#10000;
	data_in <= 24'b101010101001010001110100;
#10000;
	data_in <= 24'b101011001001100001111000;
#10000;
	data_in <= 24'b101100001001110001111011;
#10000;
	data_in <= 24'b100101101000000101100000;
#10000;
	data_in <= 24'b100110111000010101100100;
#10000;
	data_in <= 24'b100111101000100101101000;
#10000;
	data_in <= 24'b101000101000110001101100;
#10000;
	data_in <= 24'b101001011001000001110000;
#10000;
	data_in <= 24'b101010011001001101110100;
#10000;
	data_in <= 24'b101011011001011101111000;
#10000;
	data_in <= 24'b101100001001101101111011;
#10000;
	data_in <= 24'b100101101000000101100001;
#10000;
	data_in <= 24'b100110101000010101100101;
#10000;
	data_in <= 24'b100111101000100101101001;
#10000;
	data_in <= 24'b101000011000110101101101;
#10000;
	data_in <= 24'b101001011001000001110001;
#10000;
	data_in <= 24'b101010001001010001110100;
#10000;
	data_in <= 24'b101011001001011101110111;
#10000;
	data_in <= 24'b101011111001101101111011;
#10000;
	data_in <= 24'b100101101000000101100001;
#10000;
	data_in <= 24'b100110011000010001100101;
#10000;
	data_in <= 24'b100111101000100101101000;
#10000;
	data_in <= 24'b101000011000111001101100;
#10000;
	data_in <= 24'b101001001001000101110000;
#10000;
	data_in <= 24'b101001111001010101110100;
#10000;
	data_in <= 24'b101010101001100001110111;
#10000;
	data_in <= 24'b101011111001101101111011;
#10000;
	data_in <= 24'b100101101000001001011111;
#10000;
	data_in <= 24'b100110101000010101100100;
#10000;
	data_in <= 24'b100111011000100001101000;
#10000;
	data_in <= 24'b101000011000110001101011;
#10000;
	data_in <= 24'b101001001001000001101110;
#10000;
	data_in <= 24'b101001111001010001110011;
#10000;
	data_in <= 24'b101010111001011101110111;
#10000;
	data_in <= 24'b101011111001101001111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101101001001111101111111;
#10000;
	data_in <= 24'b101101101010001110000001;
#10000;
	data_in <= 24'b101110011010011010000100;
#10000;
	data_in <= 24'b101111001010100010001000;
#10000;
	data_in <= 24'b101111101010101110001011;
#10000;
	data_in <= 24'b110000101010111010001110;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b101100111001111101111111;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101110011010010110000101;
#10000;
	data_in <= 24'b101111001010100110001000;
#10000;
	data_in <= 24'b101111111010101110001011;
#10000;
	data_in <= 24'b110000101010111010001110;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b101100111001111101111110;
#10000;
	data_in <= 24'b101101101010000110000010;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101111001010100010001001;
#10000;
	data_in <= 24'b101111111010101110001011;
#10000;
	data_in <= 24'b110000011010111010001110;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110001101011001110010100;
#10000;
	data_in <= 24'b101100111001111101111110;
#10000;
	data_in <= 24'b101101101010001010000010;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101111001010011110001000;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b110000011010110110001101;
#10000;
	data_in <= 24'b110001001011000010010000;
#10000;
	data_in <= 24'b110001101011001110010100;
#10000;
	data_in <= 24'b101100111001111101111110;
#10000;
	data_in <= 24'b101101101010000110000010;
#10000;
	data_in <= 24'b101110011010010010000101;
#10000;
	data_in <= 24'b101111001010011110001000;
#10000;
	data_in <= 24'b101111101010100110001010;
#10000;
	data_in <= 24'b110000011010110010001101;
#10000;
	data_in <= 24'b110000111011000010010000;
#10000;
	data_in <= 24'b110001011011001010010011;
#10000;
	data_in <= 24'b101100101001111101111111;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101110011010010110000101;
#10000;
	data_in <= 24'b101110111010011110001000;
#10000;
	data_in <= 24'b101111101010100110001010;
#10000;
	data_in <= 24'b110000001010110110001110;
#10000;
	data_in <= 24'b110000111011000010010001;
#10000;
	data_in <= 24'b110001011011001010010011;
#10000;
	data_in <= 24'b101100101001111001111110;
#10000;
	data_in <= 24'b101101011010000110000001;
#10000;
	data_in <= 24'b101110001010010010000100;
#10000;
	data_in <= 24'b101110111010011110000111;
#10000;
	data_in <= 24'b101111011010101010001011;
#10000;
	data_in <= 24'b110000001010110110001110;
#10000;
	data_in <= 24'b110000101010111110010000;
#10000;
	data_in <= 24'b110001001011000110010010;
#10000;
	data_in <= 24'b101100101001110101111101;
#10000;
	data_in <= 24'b101101011001111101111111;
#10000;
	data_in <= 24'b101110001010001110000011;
#10000;
	data_in <= 24'b101110111010011110000111;
#10000;
	data_in <= 24'b101111011010100110001001;
#10000;
	data_in <= 24'b101111111010110010001100;
#10000;
	data_in <= 24'b110000101010111010001111;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110010001011010110010110;
#10000;
	data_in <= 24'b110010111011100010011001;
#10000;
	data_in <= 24'b110011011011101010011011;
#10000;
	data_in <= 24'b110100001011110010011101;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100101011111110100000;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b110010001011010110010110;
#10000;
	data_in <= 24'b110010111011100010011001;
#10000;
	data_in <= 24'b110011011011101110011011;
#10000;
	data_in <= 24'b110011111011110010011101;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110100111100000010100010;
#10000;
	data_in <= 24'b110101011100001010100100;
#10000;
	data_in <= 24'b110010001011010110010110;
#10000;
	data_in <= 24'b110010101011011110011000;
#10000;
	data_in <= 24'b110011001011101010011011;
#10000;
	data_in <= 24'b110011101011110010011101;
#10000;
	data_in <= 24'b110100001011111010011111;
#10000;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101011100001010100100;
#10000;
	data_in <= 24'b110010001011010110010110;
#10000;
	data_in <= 24'b110010101011011110011000;
#10000;
	data_in <= 24'b110011001011100110011010;
#10000;
	data_in <= 24'b110011011011101110011100;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100111100000010100010;
#10000;
	data_in <= 24'b110101011100001010100100;
#10000;
	data_in <= 24'b110001111011010010010101;
#10000;
	data_in <= 24'b110010011011011010011000;
#10000;
	data_in <= 24'b110010111011100010011001;
#10000;
	data_in <= 24'b110011011011101010011100;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110100101011111110100010;
#10000;
	data_in <= 24'b110101001100001010100011;
#10000;
	data_in <= 24'b110001111011010010010101;
#10000;
	data_in <= 24'b110010011011011010011000;
#10000;
	data_in <= 24'b110010111011100010011010;
#10000;
	data_in <= 24'b110011011011101010011101;
#10000;
	data_in <= 24'b110011101011110010011110;
#10000;
	data_in <= 24'b110100001011110110100000;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100101100000110100011;
#10000;
	data_in <= 24'b110001101011001110010100;
#10000;
	data_in <= 24'b110010001011011010010110;
#10000;
	data_in <= 24'b110010101011100010011010;
#10000;
	data_in <= 24'b110011001011101010011100;
#10000;
	data_in <= 24'b110011101011110010011110;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110100001011111110100000;
#10000;
	data_in <= 24'b110100101100000110100010;
#10000;
	data_in <= 24'b110001101011001110010011;
#10000;
	data_in <= 24'b110010001011010110010110;
#10000;
	data_in <= 24'b110010101011011010011000;
#10000;
	data_in <= 24'b110011001011100110011011;
#10000;
	data_in <= 24'b110011101011101110011101;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110100011011111110100000;
#10000;
	data_in <= 24'b110100101100000010100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110110101100100010101010;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111011100101110101101;
#10000;
	data_in <= 24'b110101101100001110100110;
#10000;
	data_in <= 24'b110101111100011010100111;
#10000;
	data_in <= 24'b110110011100011110101000;
#10000;
	data_in <= 24'b110110101100100010101010;
#10000;
	data_in <= 24'b110110111100100110101011;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110110001100011010100111;
#10000;
	data_in <= 24'b110110011100011010101001;
#10000;
	data_in <= 24'b110110101100011110101010;
#10000;
	data_in <= 24'b110110111100100010101011;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110101101100010010100101;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110101100011110101010;
#10000;
	data_in <= 24'b110110111100100010101011;
#10000;
	data_in <= 24'b110110111100100010101011;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100100110101101;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b110110001100010110100111;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110011100011010101000;
#10000;
	data_in <= 24'b110110101100011110101010;
#10000;
	data_in <= 24'b110110111100100010101011;
#10000;
	data_in <= 24'b110110111100100010101011;
#10000;
	data_in <= 24'b110111001100100110101101;
#10000;
	data_in <= 24'b110101001100001110100110;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110110001100010110101000;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110110101100011110101010;
#10000;
	data_in <= 24'b110110101100100010101010;
#10000;
	data_in <= 24'b110110111100100010101011;
#10000;
	data_in <= 24'b110110111100100110101100;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101111100011010101000;
#10000;
	data_in <= 24'b110110011100011110101001;
#10000;
	data_in <= 24'b110110101100100010101010;
#10000;
	data_in <= 24'b110110101100100010101011;
#10000;
	data_in <= 24'b110110111100100110101100;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101011100001110100100;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110110011100011010101010;
#10000;
	data_in <= 24'b110110011100011110101010;
#10000;
	data_in <= 24'b110110101100100010101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110111011100110010101110;
#10000;
	data_in <= 24'b110111101100110110101111;
#10000;
	data_in <= 24'b110111011100110010101111;
#10000;
	data_in <= 24'b110111111100110110101111;
#10000;
	data_in <= 24'b111000011100111010110000;
#10000;
	data_in <= 24'b101111111011110010101101;
#10000;
	data_in <= 24'b100101101010100010101011;
#10000;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110111011100110010101110;
#10000;
	data_in <= 24'b110111011100110110101111;
#10000;
	data_in <= 24'b110111111100110110101111;
#10000;
	data_in <= 24'b110111111100110110101111;
#10000;
	data_in <= 24'b101010001011000010101010;
#10000;
	data_in <= 24'b100000111001111010101011;
#10000;
	data_in <= 24'b100001111010001110101111;
#10000;
	data_in <= 24'b110111011100101110101111;
#10000;
	data_in <= 24'b110111011100110010101111;
#10000;
	data_in <= 24'b110111001100110010101111;
#10000;
	data_in <= 24'b111000011100111010110000;
#10000;
	data_in <= 24'b101011011011001010101000;
#10000;
	data_in <= 24'b011111001001101010101000;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b100011101010011110110000;
#10000;
	data_in <= 24'b110111011100101010101110;
#10000;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110111101100110110101111;
#10000;
	data_in <= 24'b110111011100110010101111;
#10000;
	data_in <= 24'b100010001001101110100000;
#10000;
	data_in <= 24'b100000001001101110100111;
#10000;
	data_in <= 24'b100011001010011010101111;
#10000;
	data_in <= 24'b100011001010010110101111;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b111000011100111010101111;
#10000;
	data_in <= 24'b100111001010010110011111;
#10000;
	data_in <= 24'b011010101000101010011010;
#10000;
	data_in <= 24'b100000001001101110100110;
#10000;
	data_in <= 24'b100001011001111110101001;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b110110111100101010101110;
#10000;
	data_in <= 24'b110111111100110010101111;
#10000;
	data_in <= 24'b110100111100010110101011;
#10000;
	data_in <= 24'b100011011001101110011010;
#10000;
	data_in <= 24'b011011011000100110010101;
#10000;
	data_in <= 24'b011010111000100110010111;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110110111100101010101101;
#10000;
	data_in <= 24'b110110111100101010101101;
#10000;
	data_in <= 24'b110111101100110010101110;
#10000;
	data_in <= 24'b110110101100101010101100;
#10000;
	data_in <= 24'b101111111011100010100100;
#10000;
	data_in <= 24'b101010101010101110011101;
#10000;
	data_in <= 24'b110110101100100110101011;
#10000;
	data_in <= 24'b110110101100100110101011;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110110101100100110101011;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b111000011100110110101110;
#10000;
	data_in <= 24'b111000001100110010101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010001010000110101100;
#10000;
	data_in <= 24'b100001111010000010101010;
#10000;
	data_in <= 24'b100000001001100010100001;
#10000;
	data_in <= 24'b100000011001011110100000;
#10000;
	data_in <= 24'b100010101001111110101001;
#10000;
	data_in <= 24'b100100111010100010110010;
#10000;
	data_in <= 24'b100110101010111010111000;
#10000;
	data_in <= 24'b100111111011001010111101;
#10000;
	data_in <= 24'b100011001010011010110000;
#10000;
	data_in <= 24'b100011011010011010101111;
#10000;
	data_in <= 24'b100010001010000010101001;
#10000;
	data_in <= 24'b100000011001100010100001;
#10000;
	data_in <= 24'b011111011001010010011101;
#10000;
	data_in <= 24'b100000001001011010011111;
#10000;
	data_in <= 24'b100001101001110010100100;
#10000;
	data_in <= 24'b100011001010000110101010;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b100011001010010110101111;
#10000;
	data_in <= 24'b100010011010000110101100;
#10000;
	data_in <= 24'b100001011001110110100110;
#10000;
	data_in <= 24'b100000011001100110100001;
#10000;
	data_in <= 24'b011111111001011010011111;
#10000;
	data_in <= 24'b011110111001010010011110;
#10000;
	data_in <= 24'b100011001010010110101111;
#10000;
	data_in <= 24'b100011001010010110101111;
#10000;
	data_in <= 24'b100010111010010110101111;
#10000;
	data_in <= 24'b100010101010010010101101;
#10000;
	data_in <= 24'b100001111010000010101001;
#10000;
	data_in <= 24'b100000001001101010100101;
#10000;
	data_in <= 24'b011101101001001010011110;
#10000;
	data_in <= 24'b011011001000100010010101;
#10000;
	data_in <= 24'b100001101001111110101001;
#10000;
	data_in <= 24'b100001011001111010101001;
#10000;
	data_in <= 24'b100000011001101110100111;
#10000;
	data_in <= 24'b011110111001011110100011;
#10000;
	data_in <= 24'b011100101001000010011101;
#10000;
	data_in <= 24'b011011001000100010010110;
#10000;
	data_in <= 24'b011011111000011010001101;
#10000;
	data_in <= 24'b100000101000101110000100;
#10000;
	data_in <= 24'b011010111000101010010111;
#10000;
	data_in <= 24'b011010111000100110010111;
#10000;
	data_in <= 24'b011010111000100010010100;
#10000;
	data_in <= 24'b011011111000100010010000;
#10000;
	data_in <= 24'b011110111000110010001101;
#10000;
	data_in <= 24'b100100101001100010001101;
#10000;
	data_in <= 24'b101011101010100010010011;
#10000;
	data_in <= 24'b101111111011010110011100;
#10000;
	data_in <= 24'b101000101010010010011010;
#10000;
	data_in <= 24'b101000111010010010011000;
#10000;
	data_in <= 24'b101010101010100110011000;
#10000;
	data_in <= 24'b101101101010111110011010;
#10000;
	data_in <= 24'b110001011011100110011111;
#10000;
	data_in <= 24'b110100011100001010100110;
#10000;
	data_in <= 24'b110101111100100010101100;
#10000;
	data_in <= 24'b110110011100100110101110;
#10000;
	data_in <= 24'b110111101100101010101100;
#10000;
	data_in <= 24'b110111011100100110101100;
#10000;
	data_in <= 24'b110111011100101010101100;
#10000;
	data_in <= 24'b110111011100101010101101;
#10000;
	data_in <= 24'b110111001100101110101111;
#10000;
	data_in <= 24'b110111001100101010101111;
#10000;
	data_in <= 24'b110111001100101010101110;
#10000;
	data_in <= 24'b110111001100101010101110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101000011011010111000000;
#10000;
	data_in <= 24'b101000101011011011000000;
#10000;
	data_in <= 24'b101000101011011011000001;
#10000;
	data_in <= 24'b101000111011011111000001;
#10000;
	data_in <= 24'b101000111011011111000001;
#10000;
	data_in <= 24'b101000101011011011000001;
#10000;
	data_in <= 24'b101000101011011011000000;
#10000;
	data_in <= 24'b101000001011010010111110;
#10000;
	data_in <= 24'b100100011010010110101110;
#10000;
	data_in <= 24'b100101011010101010110100;
#10000;
	data_in <= 24'b100110001010110110111001;
#10000;
	data_in <= 24'b100110001010110110111000;
#10000;
	data_in <= 24'b100101111010110110111000;
#10000;
	data_in <= 24'b100101101010101110110110;
#10000;
	data_in <= 24'b100100111010100010110011;
#10000;
	data_in <= 24'b100011101010001110101101;
#10000;
	data_in <= 24'b011101011001000110011101;
#10000;
	data_in <= 24'b011101001000101110010010;
#10000;
	data_in <= 24'b011110111000110010001100;
#10000;
	data_in <= 24'b011111111000111110010000;
#10000;
	data_in <= 24'b100000011001000010010000;
#10000;
	data_in <= 24'b011111101000110010001010;
#10000;
	data_in <= 24'b011101011000011110001001;
#10000;
	data_in <= 24'b011100011000110010011000;
#10000;
	data_in <= 24'b011010111000000110000100;
#10000;
	data_in <= 24'b011101100111111001110100;
#10000;
	data_in <= 24'b100000101000010101110101;
#10000;
	data_in <= 24'b100100011001000110000000;
#10000;
	data_in <= 24'b100111011001101010000110;
#10000;
	data_in <= 24'b100110011001011110000100;
#10000;
	data_in <= 24'b100010011000101001111010;
#10000;
	data_in <= 24'b011101011000001101111111;
#10000;
	data_in <= 24'b100101101001010110000011;
#10000;
	data_in <= 24'b101001001010000010001100;
#10000;
	data_in <= 24'b101100111010110010011000;
#10000;
	data_in <= 24'b110001001011100110100010;
#10000;
	data_in <= 24'b110100001100001010100111;
#10000;
	data_in <= 24'b110011111100000110100111;
#10000;
	data_in <= 24'b110000011011010110011110;
#10000;
	data_in <= 24'b101010101010001110001110;
#10000;
	data_in <= 24'b110010001011110010100011;
#10000;
	data_in <= 24'b110011111100000110101000;
#10000;
	data_in <= 24'b110101101100011010101100;
#10000;
	data_in <= 24'b110110111100101010101110;
#10000;
	data_in <= 24'b110111011100110010101111;
#10000;
	data_in <= 24'b110111011100110010101111;
#10000;
	data_in <= 24'b110111001100101010101110;
#10000;
	data_in <= 24'b110101001100010010101010;
#10000;
	data_in <= 24'b110110111100101010101110;
#10000;
	data_in <= 24'b110111001100101110101111;
#10000;
	data_in <= 24'b110111001100101110101111;
#10000;
	data_in <= 24'b110111001100101110101111;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b110111001100101010101110;
#10000;
	data_in <= 24'b110111011100101110101110;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b110111001100101110101110;
#10000;
	data_in <= 24'b110111001100101110101101;
#10000;
	data_in <= 24'b110111001100101110101101;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100111001011000010111010;
#10000;
	data_in <= 24'b100101101010101110110101;
#10000;
	data_in <= 24'b100011111010001110101110;
#10000;
	data_in <= 24'b100001001001101010100011;
#10000;
	data_in <= 24'b100000001001011010011111;
#10000;
	data_in <= 24'b100001001001110110100110;
#10000;
	data_in <= 24'b100010111010010110101110;
#10000;
	data_in <= 24'b100010001010001010101101;
#10000;
	data_in <= 24'b100010011001111010100111;
#10000;
	data_in <= 24'b100000101001100010100001;
#10000;
	data_in <= 24'b011111011001001110011100;
#10000;
	data_in <= 24'b011111011001010010011101;
#10000;
	data_in <= 24'b100001001001110010100101;
#10000;
	data_in <= 24'b100010111010010010101110;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b011101111001000110011100;
#10000;
	data_in <= 24'b011111011001010010011110;
#10000;
	data_in <= 24'b100000011001100110100010;
#10000;
	data_in <= 24'b100001101001111110101000;
#10000;
	data_in <= 24'b100010111010001110101101;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b011011011000011110010001;
#10000;
	data_in <= 24'b011100111001000010011101;
#10000;
	data_in <= 24'b011111101001100110100100;
#10000;
	data_in <= 24'b100001111010000010101010;
#10000;
	data_in <= 24'b100010111010010010101101;
#10000;
	data_in <= 24'b100011001010010110101110;
#10000;
	data_in <= 24'b100011001010010110101111;
#10000;
	data_in <= 24'b100011001010010110101111;
#10000;
	data_in <= 24'b100100101001010010000110;
#10000;
	data_in <= 24'b011111011000110110001101;
#10000;
	data_in <= 24'b011100001000101010010101;
#10000;
	data_in <= 24'b011100001000111010011100;
#10000;
	data_in <= 24'b011110001001011010100010;
#10000;
	data_in <= 24'b100000001001101110100110;
#10000;
	data_in <= 24'b100001001001111010101000;
#10000;
	data_in <= 24'b100001101010000010101001;
#10000;
	data_in <= 24'b110010011011101110100010;
#10000;
	data_in <= 24'b110000011011010110011100;
#10000;
	data_in <= 24'b101011001010100110010111;
#10000;
	data_in <= 24'b100011101001100010010010;
#10000;
	data_in <= 24'b011101111000110110010001;
#10000;
	data_in <= 24'b011011011000100110010100;
#10000;
	data_in <= 24'b011011001000100110010111;
#10000;
	data_in <= 24'b011011001000101010011000;
#10000;
	data_in <= 24'b110110101100100110101110;
#10000;
	data_in <= 24'b110110011100100010101110;
#10000;
	data_in <= 24'b110110101100100110101100;
#10000;
	data_in <= 24'b110100111100001110100110;
#10000;
	data_in <= 24'b110000101011011110011110;
#10000;
	data_in <= 24'b101011111010101110010111;
#10000;
	data_in <= 24'b101000001010001010010100;
#10000;
	data_in <= 24'b100110001001110110010010;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110110111100101010101101;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110110111100100110101010;
#10000;
	data_in <= 24'b110110011100011110101000;
#10000;
	data_in <= 24'b110101111100011010101000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011111011001101010100110;
#10000;
	data_in <= 24'b011010101000110010011100;
#10000;
	data_in <= 24'b010111111000000110010001;
#10000;
	data_in <= 24'b010111100111111110001110;
#10000;
	data_in <= 24'b010110000111101110001100;
#10000;
	data_in <= 24'b010101100111100110001011;
#10000;
	data_in <= 24'b010100100111011110001010;
#10000;
	data_in <= 24'b010011100111010010001001;
#10000;
	data_in <= 24'b100011101010011110110000;
#10000;
	data_in <= 24'b100010111010010010101101;
#10000;
	data_in <= 24'b100001001001101010100001;
#10000;
	data_in <= 24'b101011101010101010011001;
#10000;
	data_in <= 24'b110000101011010010011010;
#10000;
	data_in <= 24'b101110001010111010011000;
#10000;
	data_in <= 24'b101011111010100010010100;
#10000;
	data_in <= 24'b100111111001111010010000;
#10000;
	data_in <= 24'b100011011010011010110000;
#10000;
	data_in <= 24'b100011101010011010110000;
#10000;
	data_in <= 24'b100000011001111010101010;
#10000;
	data_in <= 24'b100010111001111010100010;
#10000;
	data_in <= 24'b110101011100010010101001;
#10000;
	data_in <= 24'b111000001100101010101011;
#10000;
	data_in <= 24'b110110111100100010101000;
#10000;
	data_in <= 24'b110110101100010110100110;
#10000;
	data_in <= 24'b100011001010010110101111;
#10000;
	data_in <= 24'b100010111010010110101110;
#10000;
	data_in <= 24'b100001111010000010101001;
#10000;
	data_in <= 24'b011011101000110010011010;
#10000;
	data_in <= 24'b101101011011000110100000;
#10000;
	data_in <= 24'b110111101100100010101001;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101101100010010100101;
#10000;
	data_in <= 24'b100001011001111110101001;
#10000;
	data_in <= 24'b100000111001110010100111;
#10000;
	data_in <= 24'b011100111001000110011111;
#10000;
	data_in <= 24'b011011101000100010010010;
#10000;
	data_in <= 24'b110000001011010110011110;
#10000;
	data_in <= 24'b110111001100100010101001;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b011010111000100110011000;
#10000;
	data_in <= 24'b011010101000011110010100;
#10000;
	data_in <= 24'b011011101000011010001111;
#10000;
	data_in <= 24'b100111111010000010010100;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110110001100011010101000;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101001100001110100110;
#10000;
	data_in <= 24'b100110011001110110010011;
#10000;
	data_in <= 24'b101001101010010110010110;
#10000;
	data_in <= 24'b101111101011010010011100;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110101101100010010100111;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110110001100011010101000;
#10000;
	data_in <= 24'b110110111100011110101010;
#10000;
	data_in <= 24'b110110111100011110101010;
#10000;
	data_in <= 24'b110110001100010110101000;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101011100001110100100;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010011100111010110001001;
#10000;
	data_in <= 24'b010110010111101010001010;
#10000;
	data_in <= 24'b011100111000100010001101;
#10000;
	data_in <= 24'b101001001010001110010101;
#10000;
	data_in <= 24'b110100011011110010011100;
#10000;
	data_in <= 24'b110100011011110010011011;
#10000;
	data_in <= 24'b110010101011100010011000;
#10000;
	data_in <= 24'b110010001011010110010110;
#10000;
	data_in <= 24'b100001011001000010001011;
#10000;
	data_in <= 24'b011001100111111110000111;
#10000;
	data_in <= 24'b010011100111001010000110;
#10000;
	data_in <= 24'b010011000111000110000110;
#10000;
	data_in <= 24'b011110101000101110001100;
#10000;
	data_in <= 24'b110001011011011010011001;
#10000;
	data_in <= 24'b110011011011101010011001;
#10000;
	data_in <= 24'b110010001011010010010110;
#10000;
	data_in <= 24'b110101011100000010100000;
#10000;
	data_in <= 24'b110001001011001110010111;
#10000;
	data_in <= 24'b100110011001100110001100;
#10000;
	data_in <= 24'b011000100111110010000110;
#10000;
	data_in <= 24'b010001100110111010000101;
#10000;
	data_in <= 24'b011101101000100010001010;
#10000;
	data_in <= 24'b110010011011011010011000;
#10000;
	data_in <= 24'b110010011011011010010110;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101101100001010100100;
#10000;
	data_in <= 24'b110101101100000010011111;
#10000;
	data_in <= 24'b101100011010011110010000;
#10000;
	data_in <= 24'b011001000111110110000110;
#10000;
	data_in <= 24'b010010100111000010000101;
#10000;
	data_in <= 24'b100111011001110010001110;
#10000;
	data_in <= 24'b110011111011100110010111;
#10000;
	data_in <= 24'b110100111100000110100011;
#10000;
	data_in <= 24'b110100001011111110100001;
#10000;
	data_in <= 24'b110011111011111010100001;
#10000;
	data_in <= 24'b110101101011111110011111;
#10000;
	data_in <= 24'b101000011001111010001100;
#10000;
	data_in <= 24'b010011110111001010000100;
#10000;
	data_in <= 24'b011100111000011010001001;
#10000;
	data_in <= 24'b110010111011010110010101;
#10000;
	data_in <= 24'b110100101100000110100011;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110011101011110010011111;
#10000;
	data_in <= 24'b110100001011110110100000;
#10000;
	data_in <= 24'b110010001011010110010111;
#10000;
	data_in <= 24'b011001110111111110000111;
#10000;
	data_in <= 24'b011000010111110010001000;
#10000;
	data_in <= 24'b110000001010111110010010;
#10000;
	data_in <= 24'b110100101100000110100010;
#10000;
	data_in <= 24'b110100001011111110100000;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110011011011110010011110;
#10000;
	data_in <= 24'b110100001011110010011011;
#10000;
	data_in <= 24'b011101101000100110001011;
#10000;
	data_in <= 24'b010110010111100110000111;
#10000;
	data_in <= 24'b101110111010110010010000;
#10000;
	data_in <= 24'b110100101100000010100010;
#10000;
	data_in <= 24'b110100011011111110100000;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110011011011101010011101;
#10000;
	data_in <= 24'b110100011011101110011011;
#10000;
	data_in <= 24'b100011011001001110001011;
#10000;
	data_in <= 24'b011100001000001010000101;
#10000;
	data_in <= 24'b110000101010111110010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110000101010111010001110;
#10000;
	data_in <= 24'b101111101010101110001011;
#10000;
	data_in <= 24'b101111001010100010001000;
#10000;
	data_in <= 24'b101110011010011010000100;
#10000;
	data_in <= 24'b101101101010001110000001;
#10000;
	data_in <= 24'b101101001001111101111111;
#10000;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110000101010111010001110;
#10000;
	data_in <= 24'b101111111010101110001011;
#10000;
	data_in <= 24'b101111001010100110001000;
#10000;
	data_in <= 24'b101110011010010110000101;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101100111001111101111111;
#10000;
	data_in <= 24'b110001101011001110010100;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110000011010111010001110;
#10000;
	data_in <= 24'b101111111010101110001011;
#10000;
	data_in <= 24'b101111001010100010001001;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101101101010000110000010;
#10000;
	data_in <= 24'b101100111001111101111110;
#10000;
	data_in <= 24'b110001001011001010010011;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110000011010110110001101;
#10000;
	data_in <= 24'b101111101010101010001010;
#10000;
	data_in <= 24'b101111001010011110001000;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101101101010001010000010;
#10000;
	data_in <= 24'b101100111001111101111110;
#10000;
	data_in <= 24'b110001011011001010010100;
#10000;
	data_in <= 24'b110000111011000010010000;
#10000;
	data_in <= 24'b110000011010110010001101;
#10000;
	data_in <= 24'b101111101010100110001010;
#10000;
	data_in <= 24'b101111001010011110001000;
#10000;
	data_in <= 24'b101110011010010010000101;
#10000;
	data_in <= 24'b101101101010000110000010;
#10000;
	data_in <= 24'b101100111001111101111110;
#10000;
	data_in <= 24'b110001111011010010010011;
#10000;
	data_in <= 24'b110000101010111110010001;
#10000;
	data_in <= 24'b110000001010110110001110;
#10000;
	data_in <= 24'b101111101010100110001010;
#10000;
	data_in <= 24'b101110111010011110001000;
#10000;
	data_in <= 24'b101110011010010110000101;
#10000;
	data_in <= 24'b101101101010001010000001;
#10000;
	data_in <= 24'b101100101001111101111111;
#10000;
	data_in <= 24'b110010001011001110010011;
#10000;
	data_in <= 24'b110000011010111010010000;
#10000;
	data_in <= 24'b110000001010110110001110;
#10000;
	data_in <= 24'b101111011010101010001011;
#10000;
	data_in <= 24'b101110111010011110000111;
#10000;
	data_in <= 24'b101110001010010010000100;
#10000;
	data_in <= 24'b101101011010000110000001;
#10000;
	data_in <= 24'b101100101001111001111110;
#10000;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b110000011010111010001111;
#10000;
	data_in <= 24'b101111111010110010001100;
#10000;
	data_in <= 24'b101111011010100110001001;
#10000;
	data_in <= 24'b101110111010011110000111;
#10000;
	data_in <= 24'b101110001010001110000011;
#10000;
	data_in <= 24'b101101011001111101111111;
#10000;
	data_in <= 24'b101100101001110101111101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101100001001101101111100;
#10000;
	data_in <= 24'b101011011001100001110111;
#10000;
	data_in <= 24'b101010101001010101110011;
#10000;
	data_in <= 24'b101001111001000101110000;
#10000;
	data_in <= 24'b101000111000110101101100;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b100110111000011001100100;
#10000;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b101100001001110001111011;
#10000;
	data_in <= 24'b101011011001100101111000;
#10000;
	data_in <= 24'b101010101001010101110100;
#10000;
	data_in <= 24'b101001111001000101110000;
#10000;
	data_in <= 24'b101000101000110101101011;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b100110111000011001100100;
#10000;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b101100001001110001111011;
#10000;
	data_in <= 24'b101011011001100101111000;
#10000;
	data_in <= 24'b101010101001010001110101;
#10000;
	data_in <= 24'b101001101001000001110001;
#10000;
	data_in <= 24'b101000101000110101101101;
#10000;
	data_in <= 24'b100111111000101001101001;
#10000;
	data_in <= 24'b100110101000010101100100;
#10000;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b101100001001110001111011;
#10000;
	data_in <= 24'b101011001001100001111000;
#10000;
	data_in <= 24'b101010101001010001110100;
#10000;
	data_in <= 24'b101001101001000101110001;
#10000;
	data_in <= 24'b101000011000110001101101;
#10000;
	data_in <= 24'b100111111000101001101000;
#10000;
	data_in <= 24'b100110101000010101100011;
#10000;
	data_in <= 24'b100101111000001001100000;
#10000;
	data_in <= 24'b101100001001101101111011;
#10000;
	data_in <= 24'b101011011001011101111000;
#10000;
	data_in <= 24'b101010011001001101110100;
#10000;
	data_in <= 24'b101001011001000001110000;
#10000;
	data_in <= 24'b101000101000110001101100;
#10000;
	data_in <= 24'b100111101000100101101000;
#10000;
	data_in <= 24'b100110111000010101100100;
#10000;
	data_in <= 24'b100101101000000101100000;
#10000;
	data_in <= 24'b101011111001101101111011;
#10000;
	data_in <= 24'b101011001001011101110111;
#10000;
	data_in <= 24'b101010001001010001110100;
#10000;
	data_in <= 24'b101001011001000001110001;
#10000;
	data_in <= 24'b101000011000110101101101;
#10000;
	data_in <= 24'b100111101000100101101001;
#10000;
	data_in <= 24'b100110101000010101100101;
#10000;
	data_in <= 24'b100101101000000101100001;
#10000;
	data_in <= 24'b101011111001101101111011;
#10000;
	data_in <= 24'b101010101001100001110111;
#10000;
	data_in <= 24'b101001111001010101110100;
#10000;
	data_in <= 24'b101001001001000101110000;
#10000;
	data_in <= 24'b101000011000111001101100;
#10000;
	data_in <= 24'b100111101000100101101000;
#10000;
	data_in <= 24'b100110011000010001100101;
#10000;
	data_in <= 24'b100101101000000101100001;
#10000;
	data_in <= 24'b101011111001101001111010;
#10000;
	data_in <= 24'b101010111001011101110111;
#10000;
	data_in <= 24'b101001111001010001110011;
#10000;
	data_in <= 24'b101001001001000001101110;
#10000;
	data_in <= 24'b101000011000110001101011;
#10000;
	data_in <= 24'b100111011000100001101000;
#10000;
	data_in <= 24'b100110101000010101100100;
#10000;
	data_in <= 24'b100101101000001001011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100101111000000101011111;
#10000;
	data_in <= 24'b100110101000010101100011;
#10000;
	data_in <= 24'b100111101000100101101000;
#10000;
	data_in <= 24'b101000011000110001101011;
#10000;
	data_in <= 24'b101001001000111101101111;
#10000;
	data_in <= 24'b101010001001010001110010;
#10000;
	data_in <= 24'b101010111001011001110110;
#10000;
	data_in <= 24'b101011101001100101111010;
#10000;
	data_in <= 24'b100101101000000101100000;
#10000;
	data_in <= 24'b100110011000010001100011;
#10000;
	data_in <= 24'b100111011000100001101000;
#10000;
	data_in <= 24'b101000001000101101101100;
#10000;
	data_in <= 24'b101001001000111001101111;
#10000;
	data_in <= 24'b101010001001001101110011;
#10000;
	data_in <= 24'b101010111001011001110110;
#10000;
	data_in <= 24'b101011101001100101111010;
#10000;
	data_in <= 24'b100101101000000001100000;
#10000;
	data_in <= 24'b100110011000001101100011;
#10000;
	data_in <= 24'b100111011000011101100111;
#10000;
	data_in <= 24'b101000011000101101101100;
#10000;
	data_in <= 24'b101001001000111001101111;
#10000;
	data_in <= 24'b101001111001000101110010;
#10000;
	data_in <= 24'b101010101001010001110101;
#10000;
	data_in <= 24'b101011011001100001111000;
#10000;
	data_in <= 24'b100101011000000001011111;
#10000;
	data_in <= 24'b100110011000001101100011;
#10000;
	data_in <= 24'b100111001000011101100110;
#10000;
	data_in <= 24'b101000001000101001101010;
#10000;
	data_in <= 24'b101000111000110101101101;
#10000;
	data_in <= 24'b101001101001000001110001;
#10000;
	data_in <= 24'b101010011001010001110101;
#10000;
	data_in <= 24'b101011001001011101111000;
#10000;
	data_in <= 24'b100101011000000001011111;
#10000;
	data_in <= 24'b100110001000001101100010;
#10000;
	data_in <= 24'b100111001000011101100101;
#10000;
	data_in <= 24'b100111111000101001101001;
#10000;
	data_in <= 24'b101000101000110101101100;
#10000;
	data_in <= 24'b101001011001000101110000;
#10000;
	data_in <= 24'b101010011001010001110100;
#10000;
	data_in <= 24'b101010111001011101110111;
#10000;
	data_in <= 24'b100101000111111001011110;
#10000;
	data_in <= 24'b100101111000001001100010;
#10000;
	data_in <= 24'b100110111000011101100110;
#10000;
	data_in <= 24'b100111101000101001101001;
#10000;
	data_in <= 24'b101000011000110101101101;
#10000;
	data_in <= 24'b101001001001000001110000;
#10000;
	data_in <= 24'b101001111001010001110100;
#10000;
	data_in <= 24'b101010101001011001110111;
#10000;
	data_in <= 24'b100100110111110101011110;
#10000;
	data_in <= 24'b100101111000000101100001;
#10000;
	data_in <= 24'b100110101000010101100101;
#10000;
	data_in <= 24'b100111011000100101101001;
#10000;
	data_in <= 24'b101000011000110101101101;
#10000;
	data_in <= 24'b101000111000111101101111;
#10000;
	data_in <= 24'b101001101001001001110010;
#10000;
	data_in <= 24'b101010101001011001110110;
#10000;
	data_in <= 24'b100100010111111001011110;
#10000;
	data_in <= 24'b100101011000000101100001;
#10000;
	data_in <= 24'b100110011000010001100100;
#10000;
	data_in <= 24'b100111001000100001101000;
#10000;
	data_in <= 24'b100111111000101101101011;
#10000;
	data_in <= 24'b101000101000111001101110;
#10000;
	data_in <= 24'b101001011001000101110001;
#10000;
	data_in <= 24'b101010001001010001110100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101100011001110001111101;
#10000;
	data_in <= 24'b101101001001111101111111;
#10000;
	data_in <= 24'b101101111010001110000011;
#10000;
	data_in <= 24'b101110101010011010000111;
#10000;
	data_in <= 24'b101111011010100110001001;
#10000;
	data_in <= 24'b101111111010101110001011;
#10000;
	data_in <= 24'b110000011010110110001110;
#10000;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b101100011001110001111101;
#10000;
	data_in <= 24'b101100111001111110000000;
#10000;
	data_in <= 24'b101101101010001010000011;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101111001010100010001001;
#10000;
	data_in <= 24'b101111111010101110001100;
#10000;
	data_in <= 24'b110000011010110110001101;
#10000;
	data_in <= 24'b110000111010111110010000;
#10000;
	data_in <= 24'b101100001001110001111100;
#10000;
	data_in <= 24'b101100111001111010000000;
#10000;
	data_in <= 24'b101101011010000110000010;
#10000;
	data_in <= 24'b101110001010010010000101;
#10000;
	data_in <= 24'b101110101010011010000111;
#10000;
	data_in <= 24'b101111011010100110001010;
#10000;
	data_in <= 24'b110000001010110010001101;
#10000;
	data_in <= 24'b110000101010111010010000;
#10000;
	data_in <= 24'b101011111001101101111011;
#10000;
	data_in <= 24'b101100101001111101111111;
#10000;
	data_in <= 24'b101101001010000010000001;
#10000;
	data_in <= 24'b101101111010001110000100;
#10000;
	data_in <= 24'b101110101010011010000111;
#10000;
	data_in <= 24'b101111001010100010001001;
#10000;
	data_in <= 24'b101111101010101010001100;
#10000;
	data_in <= 24'b110000001010110110001110;
#10000;
	data_in <= 24'b101011101001101001111010;
#10000;
	data_in <= 24'b101100001001111001111100;
#10000;
	data_in <= 24'b101100111010000001111111;
#10000;
	data_in <= 24'b101101101010001110000011;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101110111010100010001001;
#10000;
	data_in <= 24'b101111011010101010001011;
#10000;
	data_in <= 24'b101111111010110010001100;
#10000;
	data_in <= 24'b101011011001100101111010;
#10000;
	data_in <= 24'b101100001001110001111100;
#10000;
	data_in <= 24'b101100101001111101111111;
#10000;
	data_in <= 24'b101101001010001010000010;
#10000;
	data_in <= 24'b101101111010010010000101;
#10000;
	data_in <= 24'b101110101010011110001000;
#10000;
	data_in <= 24'b101111001010100110001010;
#10000;
	data_in <= 24'b101111101010101110001100;
#10000;
	data_in <= 24'b101011001001100001111000;
#10000;
	data_in <= 24'b101011101001101001111100;
#10000;
	data_in <= 24'b101100101001111001111111;
#10000;
	data_in <= 24'b101100111010000010000001;
#10000;
	data_in <= 24'b101101101010001010000100;
#10000;
	data_in <= 24'b101110001010010110000110;
#10000;
	data_in <= 24'b101110101010011110001001;
#10000;
	data_in <= 24'b101111001010101010001011;
#10000;
	data_in <= 24'b101010111001011101110111;
#10000;
	data_in <= 24'b101011011001100101111010;
#10000;
	data_in <= 24'b101100001001110001111110;
#10000;
	data_in <= 24'b101100101001111010000000;
#10000;
	data_in <= 24'b101101011010000010000011;
#10000;
	data_in <= 24'b101101111010001110000101;
#10000;
	data_in <= 24'b101110011010011110000111;
#10000;
	data_in <= 24'b101110111010100110001001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b110010001011010010010110;
#10000;
	data_in <= 24'b110010101011011010011000;
#10000;
	data_in <= 24'b110011001011011110011010;
#10000;
	data_in <= 24'b110011101011100110011100;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110100001011111010011111;
#10000;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110001011011000110010011;
#10000;
	data_in <= 24'b110001111011001110010101;
#10000;
	data_in <= 24'b110010001011010010010111;
#10000;
	data_in <= 24'b110010111011011010011001;
#10000;
	data_in <= 24'b110011001011100110011100;
#10000;
	data_in <= 24'b110011011011101010011101;
#10000;
	data_in <= 24'b110100001011110010011111;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110001001011000010010010;
#10000;
	data_in <= 24'b110001101011001010010100;
#10000;
	data_in <= 24'b110010001011010010010110;
#10000;
	data_in <= 24'b110010011011011010010111;
#10000;
	data_in <= 24'b110010111011100010011001;
#10000;
	data_in <= 24'b110011011011101010011100;
#10000;
	data_in <= 24'b110011111011101110011111;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110000111010111110010001;
#10000;
	data_in <= 24'b110001011011000110010011;
#10000;
	data_in <= 24'b110001111011001110010101;
#10000;
	data_in <= 24'b110010001011011010010110;
#10000;
	data_in <= 24'b110010101011011110011000;
#10000;
	data_in <= 24'b110011011011100110011011;
#10000;
	data_in <= 24'b110011101011101110011101;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110000011010111010001111;
#10000;
	data_in <= 24'b110000111011000010010001;
#10000;
	data_in <= 24'b110001011011001010010011;
#10000;
	data_in <= 24'b110001111011010010010101;
#10000;
	data_in <= 24'b110010101011011010011000;
#10000;
	data_in <= 24'b110010111011100010011001;
#10000;
	data_in <= 24'b110011011011101010011010;
#10000;
	data_in <= 24'b110011101011101110011100;
#10000;
	data_in <= 24'b101111111010110110001110;
#10000;
	data_in <= 24'b110000011011000010010000;
#10000;
	data_in <= 24'b110001001011000110010010;
#10000;
	data_in <= 24'b110001111011001110010101;
#10000;
	data_in <= 24'b110010011011010110010111;
#10000;
	data_in <= 24'b110010101011011010011001;
#10000;
	data_in <= 24'b110010111011100010011010;
#10000;
	data_in <= 24'b110011011011101010011100;
#10000;
	data_in <= 24'b101111101010110010001101;
#10000;
	data_in <= 24'b110000011010111010010000;
#10000;
	data_in <= 24'b110000111011000010010010;
#10000;
	data_in <= 24'b110001011011001010010100;
#10000;
	data_in <= 24'b110001101011001110010101;
#10000;
	data_in <= 24'b110010001011010110010111;
#10000;
	data_in <= 24'b110010011011011010011001;
#10000;
	data_in <= 24'b110010111011011110011010;
#10000;
	data_in <= 24'b101111011010101110001100;
#10000;
	data_in <= 24'b110000001010110110001111;
#10000;
	data_in <= 24'b110000011010111010010000;
#10000;
	data_in <= 24'b110000111011000010010010;
#10000;
	data_in <= 24'b110001011011001010010100;
#10000;
	data_in <= 24'b110001101011001110010101;
#10000;
	data_in <= 24'b110001111011010010010110;
#10000;
	data_in <= 24'b110010001011010110010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101001100000110100100;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110110001100010110101000;
#10000;
	data_in <= 24'b110110001100011010101010;
#10000;
	data_in <= 24'b110110011100011110101010;
#10000;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101001100000110100100;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101111100010010101000;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110100101011111010100001;
#10000;
	data_in <= 24'b110101001100000010100011;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101101100001110100111;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110100001011110110011111;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110100101011111010100001;
#10000;
	data_in <= 24'b110100111011111110100011;
#10000;
	data_in <= 24'b110100111100000010100011;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110011111011110010011101;
#10000;
	data_in <= 24'b110100001011110110011111;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110100111100000010100011;
#10000;
	data_in <= 24'b110100111100000110100011;
#10000;
	data_in <= 24'b110100111100000110100011;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110011101011101110011101;
#10000;
	data_in <= 24'b110011111011110010011101;
#10000;
	data_in <= 24'b110100001011110110011111;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100101100000010100010;
#10000;
	data_in <= 24'b110100101100000010100011;
#10000;
	data_in <= 24'b110100111100000110100011;
#10000;
	data_in <= 24'b110011001011100010011011;
#10000;
	data_in <= 24'b110011011011100110011101;
#10000;
	data_in <= 24'b110011101011101110011110;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110010101011011010011001;
#10000;
	data_in <= 24'b110010111011100010011010;
#10000;
	data_in <= 24'b110011011011100110011101;
#10000;
	data_in <= 24'b110011011011101110011101;
#10000;
	data_in <= 24'b110011101011101110011110;
#10000;
	data_in <= 24'b110011111011110010011111;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110110011100100010101011;
#10000;
	data_in <= 24'b110110101100100010101011;
#10000;
	data_in <= 24'b110110011100100010101011;
#10000;
	data_in <= 24'b110110011100100010101011;
#10000;
	data_in <= 24'b110110011100100110101011;
#10000;
	data_in <= 24'b110110011100100010101100;
#10000;
	data_in <= 24'b110110011100100010101100;
#10000;
	data_in <= 24'b110110111100100010101100;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101010;
#10000;
	data_in <= 24'b110110011100011110101010;
#10000;
	data_in <= 24'b110110011100011110101010;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110101100011110101100;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101010;
#10000;
	data_in <= 24'b110110011100011010101010;
#10000;
	data_in <= 24'b110110011100011010101010;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110101101100010110101000;
#10000;
	data_in <= 24'b110101111100010110101001;
#10000;
	data_in <= 24'b110110001100010110101001;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110101001100001110100100;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100010010100101;
#10000;
	data_in <= 24'b110101011100010010100110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110100111100000110100100;
#10000;
	data_in <= 24'b110100111100000110100100;
#10000;
	data_in <= 24'b110100111100000110100100;
#10000;
	data_in <= 24'b110100111100000110100101;
#10000;
	data_in <= 24'b110101001100001010100101;
#10000;
	data_in <= 24'b110101001100001010100101;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110100101100000010100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100011;
#10000;
	data_in <= 24'b110100011011111110100100;
#10000;
	data_in <= 24'b110100101011111110100100;
#10000;
	data_in <= 24'b110100101011111110100100;
#10000;
	data_in <= 24'b110100101011111110100100;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110100001011111010100001;
#10000;
	data_in <= 24'b110100001011111010100001;
#10000;
	data_in <= 24'b110100001011111010100001;
#10000;
	data_in <= 24'b110100011011111010100001;
#10000;
	data_in <= 24'b110100011011111010100001;
#10000;
	data_in <= 24'b110100011011111010100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110110111100100010101100;
#10000;
	data_in <= 24'b110110111100100110101100;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110110111100101010101100;
#10000;
	data_in <= 24'b110110111100101010101101;
#10000;
	data_in <= 24'b110110111100101010101101;
#10000;
	data_in <= 24'b110110111100101010101101;
#10000;
	data_in <= 24'b110110111100101010101101;
#10000;
	data_in <= 24'b110110101100011110101100;
#10000;
	data_in <= 24'b110110101100100010101100;
#10000;
	data_in <= 24'b110110101100100010101100;
#10000;
	data_in <= 24'b110110101100100010101101;
#10000;
	data_in <= 24'b110110101100100010101101;
#10000;
	data_in <= 24'b110110101100100010101101;
#10000;
	data_in <= 24'b110110101100100010101101;
#10000;
	data_in <= 24'b110110101100100110101101;
#10000;
	data_in <= 24'b110110011100011010101010;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110101111100010110101001;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101000;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101010;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101101100010110100110;
#10000;
	data_in <= 24'b110101101100010110100110;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101101100010110101000;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110100101100000010100100;
#10000;
	data_in <= 24'b110100101100000110100011;
#10000;
	data_in <= 24'b110100101100000010100100;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101010101101;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111001100101010101100;
#10000;
	data_in <= 24'b110111001100100110101100;
#10000;
	data_in <= 24'b110111001100100010101100;
#10000;
	data_in <= 24'b110110101100100110101101;
#10000;
	data_in <= 24'b110110101100100110101101;
#10000;
	data_in <= 24'b110110101100100110101101;
#10000;
	data_in <= 24'b110110101100100110101101;
#10000;
	data_in <= 24'b110110101100100110101101;
#10000;
	data_in <= 24'b110110101100100110101100;
#10000;
	data_in <= 24'b110110101100100010101100;
#10000;
	data_in <= 24'b110110101100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011010101010;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101010;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100011010101000;
#10000;
	data_in <= 24'b110101111100011010101001;
#10000;
	data_in <= 24'b110101111100010110101001;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101101100010110101000;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101101100010110100110;
#10000;
	data_in <= 24'b110101101100010110100110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100101;
#10000;
	data_in <= 24'b110100101100000010100100;
#10000;
	data_in <= 24'b110100101100000110100011;
#10000;
	data_in <= 24'b110100101100000010100100;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110110111100100010101100;
#10000;
	data_in <= 24'b110110101100100010101100;
#10000;
	data_in <= 24'b110110101100100010101100;
#10000;
	data_in <= 24'b110110011100100010101011;
#10000;
	data_in <= 24'b110110011100100010101011;
#10000;
	data_in <= 24'b110110011100100010101011;
#10000;
	data_in <= 24'b110110101100100010101100;
#10000;
	data_in <= 24'b110110011100100010101011;
#10000;
	data_in <= 24'b110110101100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101100;
#10000;
	data_in <= 24'b110110011100011110101011;
#10000;
	data_in <= 24'b110110011100011110101010;
#10000;
	data_in <= 24'b110110011100011110101010;
#10000;
	data_in <= 24'b110110001100011010101010;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110011100011010101010;
#10000;
	data_in <= 24'b110110011100011010101010;
#10000;
	data_in <= 24'b110110001100011010101010;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110110001100010110101001;
#10000;
	data_in <= 24'b110101111100010110101001;
#10000;
	data_in <= 24'b110101101100010110101000;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110101101100010110100111;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110101111100010110100111;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101101100010010100110;
#10000;
	data_in <= 24'b110101011100010010100110;
#10000;
	data_in <= 24'b110101011100010010100101;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101001100001110100100;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101001100001010100101;
#10000;
	data_in <= 24'b110101001100001010100101;
#10000;
	data_in <= 24'b110100111100000110100101;
#10000;
	data_in <= 24'b110100111100000110100100;
#10000;
	data_in <= 24'b110100111100000110100100;
#10000;
	data_in <= 24'b110100111100000110100100;
#10000;
	data_in <= 24'b110100101011111110100100;
#10000;
	data_in <= 24'b110100101011111110100100;
#10000;
	data_in <= 24'b110100101011111110100100;
#10000;
	data_in <= 24'b110100011011111110100100;
#10000;
	data_in <= 24'b110100011011111110100011;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100011011111110100010;
#10000;
	data_in <= 24'b110100101100000010100010;
#10000;
	data_in <= 24'b110100011011111010100001;
#10000;
	data_in <= 24'b110100011011111010100001;
#10000;
	data_in <= 24'b110100011011111010100001;
#10000;
	data_in <= 24'b110100001011111010100001;
#10000;
	data_in <= 24'b110100001011111010100001;
#10000;
	data_in <= 24'b110100001011111010100001;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110110011100011110101010;
#10000;
	data_in <= 24'b110110001100011010101010;
#10000;
	data_in <= 24'b110110001100010110101000;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101111100010010100110;
#10000;
	data_in <= 24'b110101101100001110100101;
#10000;
	data_in <= 24'b110101001100000110100100;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110110001100011010101001;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110101111100010010101000;
#10000;
	data_in <= 24'b110101111100010010100111;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101001100000110100100;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110101111100010110101000;
#10000;
	data_in <= 24'b110101101100001110100111;
#10000;
	data_in <= 24'b110101011100001010100101;
#10000;
	data_in <= 24'b110101001100000110100011;
#10000;
	data_in <= 24'b110101001100000010100011;
#10000;
	data_in <= 24'b110100101011111010100001;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110101011100001110100110;
#10000;
	data_in <= 24'b110101011100001110100101;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110100111100000010100011;
#10000;
	data_in <= 24'b110100111011111110100011;
#10000;
	data_in <= 24'b110100101011111010100001;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110100001011110110011111;
#10000;
	data_in <= 24'b110101001100001010100100;
#10000;
	data_in <= 24'b110100111100000110100011;
#10000;
	data_in <= 24'b110100111100000110100011;
#10000;
	data_in <= 24'b110100111100000010100011;
#10000;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110100011011111010011111;
#10000;
	data_in <= 24'b110100001011110110011111;
#10000;
	data_in <= 24'b110011111011110010011101;
#10000;
	data_in <= 24'b110100111100000110100011;
#10000;
	data_in <= 24'b110100101100000010100011;
#10000;
	data_in <= 24'b110100101100000010100010;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110100001011110110011111;
#10000;
	data_in <= 24'b110011111011110010011101;
#10000;
	data_in <= 24'b110011101011101110011101;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100011011111110100001;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110011101011101110011110;
#10000;
	data_in <= 24'b110011011011100110011101;
#10000;
	data_in <= 24'b110011001011100010011011;
#10000;
	data_in <= 24'b110100001011111010100000;
#10000;
	data_in <= 24'b110011111011110110011111;
#10000;
	data_in <= 24'b110011111011110010011111;
#10000;
	data_in <= 24'b110011101011101110011110;
#10000;
	data_in <= 24'b110011011011101110011101;
#10000;
	data_in <= 24'b110011011011100110011101;
#10000;
	data_in <= 24'b110010111011100010011010;
#10000;
	data_in <= 24'b110010101011011010011001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110100101011111110100001;
#10000;
	data_in <= 24'b110100001011111010011111;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110011011011100110011100;
#10000;
	data_in <= 24'b110011011011100010011010;
#10000;
	data_in <= 24'b110000011010111110010010;
#10000;
	data_in <= 24'b101110011010100010001101;
#10000;
	data_in <= 24'b110001101011001010010011;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110100001011110010011111;
#10000;
	data_in <= 24'b110011011011101010011101;
#10000;
	data_in <= 24'b110011001011100110011100;
#10000;
	data_in <= 24'b110010101011011010011001;
#10000;
	data_in <= 24'b110010101011011010011000;
#10000;
	data_in <= 24'b110010011011010110010110;
#10000;
	data_in <= 24'b110001011011000110010011;
#10000;
	data_in <= 24'b110100011011110110100000;
#10000;
	data_in <= 24'b110011111011101110011111;
#10000;
	data_in <= 24'b110011011011101010011100;
#10000;
	data_in <= 24'b110010111011100010011001;
#10000;
	data_in <= 24'b110010011011011010010111;
#10000;
	data_in <= 24'b110010001011010010010110;
#10000;
	data_in <= 24'b110001011011000110010100;
#10000;
	data_in <= 24'b110001001011000010010010;
#10000;
	data_in <= 24'b110011111011110010011110;
#10000;
	data_in <= 24'b110011101011101110011101;
#10000;
	data_in <= 24'b110011011011100110011011;
#10000;
	data_in <= 24'b110010101011011110011000;
#10000;
	data_in <= 24'b110010001011011010010110;
#10000;
	data_in <= 24'b110001111011001110010101;
#10000;
	data_in <= 24'b110001011011000110010011;
#10000;
	data_in <= 24'b110000111010111110010001;
#10000;
	data_in <= 24'b110011101011101110011100;
#10000;
	data_in <= 24'b110011011011101010011010;
#10000;
	data_in <= 24'b110010111011100010011001;
#10000;
	data_in <= 24'b110010101011011010011000;
#10000;
	data_in <= 24'b110001111011010010010101;
#10000;
	data_in <= 24'b110001011011001010010011;
#10000;
	data_in <= 24'b110000111011000010010001;
#10000;
	data_in <= 24'b110000011010111010001111;
#10000;
	data_in <= 24'b110011011011101010011100;
#10000;
	data_in <= 24'b110010111011100010011010;
#10000;
	data_in <= 24'b110010101011011010011001;
#10000;
	data_in <= 24'b110010011011010110010111;
#10000;
	data_in <= 24'b110001111011001110010101;
#10000;
	data_in <= 24'b110001001011000110010010;
#10000;
	data_in <= 24'b110000011011000010010000;
#10000;
	data_in <= 24'b101111111010110110001110;
#10000;
	data_in <= 24'b110010111011011110011010;
#10000;
	data_in <= 24'b110010011011011010011001;
#10000;
	data_in <= 24'b110010001011010110010111;
#10000;
	data_in <= 24'b110001101011001110010101;
#10000;
	data_in <= 24'b110001011011001010010100;
#10000;
	data_in <= 24'b110000111011000010010010;
#10000;
	data_in <= 24'b110000011010111010010000;
#10000;
	data_in <= 24'b101111101010110010001101;
#10000;
	data_in <= 24'b110010001011010110010111;
#10000;
	data_in <= 24'b110001111011010010010110;
#10000;
	data_in <= 24'b110001101011001110010101;
#10000;
	data_in <= 24'b110001011011001010010100;
#10000;
	data_in <= 24'b110000111011000010010010;
#10000;
	data_in <= 24'b110000011010111010010000;
#10000;
	data_in <= 24'b110000001010110110001111;
#10000;
	data_in <= 24'b101111011010101110001100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110001001011000010010001;
#10000;
	data_in <= 24'b110000011010110110001110;
#10000;
	data_in <= 24'b101111111010101110001011;
#10000;
	data_in <= 24'b101111011010100110001001;
#10000;
	data_in <= 24'b101110101010011010000111;
#10000;
	data_in <= 24'b101101111010001110000011;
#10000;
	data_in <= 24'b101101001001111101111111;
#10000;
	data_in <= 24'b101100011001110001111101;
#10000;
	data_in <= 24'b110000111010111110010000;
#10000;
	data_in <= 24'b110000011010110110001110;
#10000;
	data_in <= 24'b101111111010101110001100;
#10000;
	data_in <= 24'b101111001010100010001001;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101101101010001010000011;
#10000;
	data_in <= 24'b101100111001111110000000;
#10000;
	data_in <= 24'b101100011001110001111101;
#10000;
	data_in <= 24'b110000101010111010010000;
#10000;
	data_in <= 24'b110000001010110010001101;
#10000;
	data_in <= 24'b101111011010100110001010;
#10000;
	data_in <= 24'b101110101010011010000111;
#10000;
	data_in <= 24'b101110001010010010000101;
#10000;
	data_in <= 24'b101101011010000110000010;
#10000;
	data_in <= 24'b101100111001111010000000;
#10000;
	data_in <= 24'b101100001001110001111100;
#10000;
	data_in <= 24'b110000001010110110001110;
#10000;
	data_in <= 24'b101111101010101010001100;
#10000;
	data_in <= 24'b101111001010100010001001;
#10000;
	data_in <= 24'b101110101010011010000111;
#10000;
	data_in <= 24'b101101111010001110000100;
#10000;
	data_in <= 24'b101101001010000010000001;
#10000;
	data_in <= 24'b101100101001111101111111;
#10000;
	data_in <= 24'b101011111001101101111011;
#10000;
	data_in <= 24'b101111111010110010001100;
#10000;
	data_in <= 24'b101111011010101010001011;
#10000;
	data_in <= 24'b101110111010100010001001;
#10000;
	data_in <= 24'b101110011010010110000110;
#10000;
	data_in <= 24'b101101101010001110000011;
#10000;
	data_in <= 24'b101100111010000001111111;
#10000;
	data_in <= 24'b101100001001111001111100;
#10000;
	data_in <= 24'b101011101001101001111010;
#10000;
	data_in <= 24'b101111101010101110001100;
#10000;
	data_in <= 24'b101111001010100110001010;
#10000;
	data_in <= 24'b101110101010011110001000;
#10000;
	data_in <= 24'b101101111010010010000101;
#10000;
	data_in <= 24'b101101001010001010000010;
#10000;
	data_in <= 24'b101100101001111101111111;
#10000;
	data_in <= 24'b101100001001110001111100;
#10000;
	data_in <= 24'b101011011001100101111010;
#10000;
	data_in <= 24'b101111001010101010001011;
#10000;
	data_in <= 24'b101110101010011110001001;
#10000;
	data_in <= 24'b101110001010010110000110;
#10000;
	data_in <= 24'b101101101010001010000100;
#10000;
	data_in <= 24'b101100111010000010000001;
#10000;
	data_in <= 24'b101100101001111001111111;
#10000;
	data_in <= 24'b101011101001101001111100;
#10000;
	data_in <= 24'b101011001001100001111000;
#10000;
	data_in <= 24'b101110111010100110001001;
#10000;
	data_in <= 24'b101110011010011110000111;
#10000;
	data_in <= 24'b101101111010001110000101;
#10000;
	data_in <= 24'b101101011010000010000011;
#10000;
	data_in <= 24'b101100101001111010000000;
#10000;
	data_in <= 24'b101100001001110001111110;
#10000;
	data_in <= 24'b101011011001100101111010;
#10000;
	data_in <= 24'b101010111001011101110111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
end_of_file_signal <= 1'b1;
	data_in <= 24'b101011101001100101111010;
#10000;
	data_in <= 24'b101010111001011001110110;
#10000;
	data_in <= 24'b101010001001010001110010;
#10000;
	data_in <= 24'b101001001000111101101111;
#10000;
	data_in <= 24'b101000011000110001101011;
#10000;
	data_in <= 24'b100111101000100101101000;
#10000;
	data_in <= 24'b100110101000010101100011;
#10000;
	data_in <= 24'b100101111000000101011111;
#10000;
	data_in <= 24'b101011101001100101111010;
#10000;
	data_in <= 24'b101010111001011001110110;
#10000;
	data_in <= 24'b101010001001001101110011;
#10000;
	data_in <= 24'b101001001000111001101111;
#10000;
	data_in <= 24'b101000001000101101101100;
#10000;
	data_in <= 24'b100111011000100001101000;
#10000;
	data_in <= 24'b100110011000010001100011;
#10000;
	data_in <= 24'b100101101000000101100000;
#10000;
	data_in <= 24'b101011011001100001111000;
#10000;
	data_in <= 24'b101010101001010001110101;
#10000;
	data_in <= 24'b101001111001000101110010;
#10000;
	data_in <= 24'b101001001000111001101111;
#10000;
	data_in <= 24'b101000011000101101101100;
#10000;
	data_in <= 24'b100111011000011101100111;
#10000;
	data_in <= 24'b100110011000001101100011;
#10000;
	data_in <= 24'b100101101000000001100000;
#10000;
	data_in <= 24'b101011001001011101111000;
#10000;
	data_in <= 24'b101010011001010001110101;
#10000;
	data_in <= 24'b101001101001000001110001;
#10000;
	data_in <= 24'b101000111000110101101101;
#10000;
	data_in <= 24'b101000001000101001101010;
#10000;
	data_in <= 24'b100111001000011101100110;
#10000;
	data_in <= 24'b100110011000001101100011;
#10000;
	data_in <= 24'b100101011000000001011111;
#10000;
	data_in <= 24'b101010111001011101110111;
#10000;
	data_in <= 24'b101010011001010001110100;
#10000;
	data_in <= 24'b101001011001000101110000;
#10000;
	data_in <= 24'b101000101000110101101100;
#10000;
	data_in <= 24'b100111111000101001101001;
#10000;
	data_in <= 24'b100111001000011101100101;
#10000;
	data_in <= 24'b100110001000001101100010;
#10000;
	data_in <= 24'b100101011000000001011111;
#10000;
	data_in <= 24'b101010101001011001110111;
#10000;
	data_in <= 24'b101001111001010001110100;
#10000;
	data_in <= 24'b101001001001000001110000;
#10000;
	data_in <= 24'b101000011000110101101101;
#10000;
	data_in <= 24'b100111101000101001101001;
#10000;
	data_in <= 24'b100110111000011101100110;
#10000;
	data_in <= 24'b100101111000001001100010;
#10000;
	data_in <= 24'b100101000111111001011110;
#10000;
	data_in <= 24'b101010101001011001110110;
#10000;
	data_in <= 24'b101001101001001001110010;
#10000;
	data_in <= 24'b101000111000111101101111;
#10000;
	data_in <= 24'b101000011000110101101101;
#10000;
	data_in <= 24'b100111011000100101101001;
#10000;
	data_in <= 24'b100110101000010101100101;
#10000;
	data_in <= 24'b100101111000000101100001;
#10000;
	data_in <= 24'b100100110111110101011110;
#10000;
	data_in <= 24'b101010001001010001110100;
#10000;
	data_in <= 24'b101001011001000101110001;
#10000;
	data_in <= 24'b101000101000111001101110;
#10000;
	data_in <= 24'b100111111000101101101011;
#10000;
	data_in <= 24'b100111001000100001101000;
#10000;
	data_in <= 24'b100110011000010001100100;
#10000;
	data_in <= 24'b100101011000000101100001;
#10000;
	data_in <= 24'b100100010111111001011110;
#10000;




                #130000;
        enable = 1'b0;

        #2000000;
		   yes = 1'b1;
    end

    // ----------------------
    // Open output file once
    // ----------------------
    initial begin
        outfile = $fopen("bitstream_output.txt", "w");
        if (outfile == 0) begin
            $display("ERROR: Could not open bitstream_output.txt");
            $finish;
        end
    end

    // ----------------------
    // End simulation when JPEG bitstream = 0
    // ----------------------
    always_ff @(posedge clk) begin
        if (data_ready) begin
            if (   yes == 1'b1) begin
                $display("INFO: End of JPEG stream detected. Closing file and stopping.");
                $fclose(outfile);
                $finish;
            end
        end
    end

    // ----------------------
    // Clock generator
    // ----------------------
    always begin : CLOCK_clk
        clk = 1'b0;
        #5000;
        clk = 1'b1;
        #5000;
    end

    // ----------------------
    // Write JPEG bitstream whenever ready
    // ----------------------
    always_ff @(posedge clk) begin : JPEG
        if (data_ready) begin
            $fwrite(outfile, "%h\n", JPEG_bitstream);   // write in hex
        end
    end

endmodule
