// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
//    Header file defining localparams for JPEG Huffman encoding.
//    - DC Huffman code lengths and codes (Luma & Chroma)
//    - AC Huffman code lengths and codes (Luma & Chroma)
//    - Run-length/size to Huffman index mapping
//
// Author: Rameen
// Date  : 23rd July 2025

`ifndef CB_HUFF_CONSTANTS_SVH
`define CB_HUFF_CONSTANTS_SVH

/* These Y DC and AC code lengths, run lengths, and bit codes
were created from the Huffman table entries in the JPEG file header.
For different Huffman tables for different images, these values
below will need to be changed.  I created a matlab file to automatically
create these entries from the already encoded JPEG image. This matlab program
won't be any help if you're starting from scratch with a .tif or other
raw image file format.  The values below come from a Huffman table, they
do not actually create the Huffman table based on the probabilities of
each code created from the image data.  You will need another program to
create the optimal Huffman table, or you can go with a generic Huffman table,
which will have slightly less than the best compression.*/


// For DC lengths
logic [3:0] Cb_DC_code_length [0:11] = '{2,2,2,3,4,5,6,7,8,9,10,11};

// For DC codes
logic [10:0] Cb_DC [0:11] = '{
    11'b00000000000,
    11'b01000000000,
    11'b10000000000,
    11'b11000000000,
    11'b11100000000,
    11'b11110000000,
    11'b11111000000,
    11'b11111100000,
    11'b11111110000,
    11'b11111111000,
    11'b11111111100,
    11'b11111111110
} ;

logic [4:0] Cb_AC_code_length [0:161] = '{
2 ,
2 ,
3 ,
4 ,
4 ,
4 ,
5 ,
5 ,
5 ,
6 ,
 6 ,
 7 ,
 7 ,
 7 ,
 7 ,
 8 ,
 8 ,
 8 ,
 9 ,
 9 ,
 9 ,
 9 ,
 9 ,
 10 ,
 10 ,
 10 ,
 10 ,
 10 ,
 11 ,
 11 ,
 11 ,
 11 ,
 12 ,
 12 ,
12 ,
12 ,
15 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16 ,
 16
};

logic [15:0] Cb_AC [0:161] = '{
    // First unique values
16'b0000000000000000 ,
16'b0100000000000000 ,
16'b1000000000000000 ,
16'b1010000000000000 ,
16'b1011000000000000 ,
16'b1100000000000000 ,
16'b1101000000000000 ,
16'b1101100000000000 ,
16'b1110000000000000 ,
16'b1110100000000000 ,
16'b1110110000000000 ,
16'b1111000000000000 ,
16'b1111001000000000 ,
16'b1111010000000000 ,
16'b1111011000000000 ,
16'b1111100000000000 ,
16'b1111100100000000 ,
16'b1111101000000000 ,
16'b1111101100000000 ,
16'b1111101110000000 ,
16'b1111110000000000 ,
16'b1111110010000000 ,
16'b1111110100000000 ,
16'b1111110110000000 ,
16'b1111110111000000 ,
16'b1111111000000000 ,
16'b1111111001000000 ,
16'b1111111010000000 ,
16'b1111111011000000 ,
16'b1111111011100000 ,
16'b1111111100000000 ,
16'b1111111100100000 ,
16'b1111111101000000 ,
16'b1111111101010000 ,
16'b1111111101100000 ,
16'b1111111101110000 ,
16'b1111111110000000 ,
16'b1111111110000010 ,
16'b1111111110000011 ,
16'b1111111110000100 ,
16'b1111111110000101 ,
16'b1111111110000110 ,
16'b1111111110000111 ,
16'b1111111110001000 ,
16'b1111111110001001 ,
16'b1111111110001010 ,
16'b1111111110001011 ,
16'b1111111110001100 ,
16'b1111111110001101 ,
16'b1111111110001110 ,
16'b1111111110001111 ,
16'b1111111110010000 ,
16'b1111111110010001 ,
16'b1111111110010010 ,
16'b1111111110010011 ,
16'b1111111110010100 ,
16'b1111111110010101 ,
16'b1111111110010110 ,
16'b1111111110010111 ,
16'b1111111110011000 ,
16'b1111111110011001 ,
16'b1111111110011010 ,
16'b1111111110011011 ,
16'b1111111110011100 ,
16'b1111111110011101 ,
16'b1111111110011110 ,
16'b1111111110011111 ,
16'b1111111110100000 ,
16'b1111111110100001 ,
16'b1111111110100010 ,
16'b1111111110100011 ,
16'b1111111110100100 ,
16'b1111111110100101 ,
16'b1111111110100110 ,
16'b1111111110100111 ,
16'b1111111110101000 ,
16'b1111111110101001 ,
16'b1111111110101010 ,
16'b1111111110101011 ,
16'b1111111110101100 ,
16'b1111111110101101 ,
16'b1111111110101110 ,
16'b1111111110101111 ,
16'b1111111110110000 ,
16'b1111111110110001 ,
16'b1111111110110010 ,
16'b1111111110110011 ,
16'b1111111110110100 ,
16'b1111111110110101 ,
16'b1111111110110110 ,
16'b1111111110110111 ,
16'b1111111110111000 ,
16'b1111111110111001 ,
16'b1111111110111010 ,
16'b1111111110111011 ,
16'b1111111110111100 ,
16'b1111111110111101 ,
16'b1111111110111110 ,
16'b1111111110111111 ,
16'b1111111111000000 ,
 16'b1111111111000001 ,
 16'b1111111111000010 ,
 16'b1111111111000011 ,
 16'b1111111111000100 ,
 16'b1111111111000101 ,
 16'b1111111111000110 ,
 16'b1111111111000111 ,
 16'b1111111111001000 ,
 16'b1111111111001001 ,
 16'b1111111111001010 ,
 16'b1111111111001011 ,
 16'b1111111111001100 ,
 16'b1111111111001101 ,
 16'b1111111111001110 ,
 16'b1111111111001111 ,
 16'b1111111111010000 ,
 16'b1111111111010001 ,
 16'b1111111111010010 ,
 16'b1111111111010011 ,
 16'b1111111111010100 ,
 16'b1111111111010101 ,
 16'b1111111111010110 ,
 16'b1111111111010111 ,
 16'b1111111111011000 ,
 16'b1111111111011001 ,
 16'b1111111111011010 ,
 16'b1111111111011011 ,
 16'b1111111111011100 ,
 16'b1111111111011101 ,
 16'b1111111111011110 ,
 16'b1111111111011111 ,
 16'b1111111111100000 ,
 16'b1111111111100001 ,
 16'b1111111111100010 ,
 16'b1111111111100011 ,
 16'b1111111111100100 ,
 16'b1111111111100101 ,
 16'b1111111111100110 ,
 16'b1111111111100111 ,
 16'b1111111111101000 ,
 16'b1111111111101001 ,
 16'b1111111111101010 ,
 16'b1111111111101011 ,
 16'b1111111111101100 ,
 16'b1111111111101101 ,
 16'b1111111111101110 ,
 16'b1111111111101111 ,
 16'b1111111111110000 ,
 16'b1111111111110001 ,
 16'b1111111111110010 ,
 16'b1111111111110011 ,
 16'b1111111111110100 ,
 16'b1111111111110101 ,
 16'b1111111111110110 ,
 16'b1111111111110111 ,
 16'b1111111111111000 ,
 16'b1111111111111001 ,
 16'b1111111111111010 ,
 16'b1111111111111011 ,
 16'b1111111111111100 ,
 16'b1111111111111101 ,
 16'b1111111111111110
};

// Define Cb_AC_run_code as a constant arraCb
localparam logic [7:0] Cb_AC_run_code [0:250] = '{
    8'd3,   // [0]
    8'd0,   // [1]
    8'd1,   // [2]
    8'd2,   // [3]
    8'd4,   // [4]
    8'd6,   // [5]
    8'd11,  // [6]
    8'd15,  // [7]
    8'd23,  // [8]
    8'd37,  // [9]
    8'd38,  // [10]
    8'd0,   // [11]
    8'd0,   // [12]
    8'd0,   // [13]
    8'd0,   // [14]
    8'd0,   // [15]
    8'd0,   // [16]
    8'd5,   // [17]
    8'd7,   // [18]
    8'd12,  // [19]
    8'd18,  // [20]
    8'd28,  // [21]
    8'd39,  // [22]
    8'd40,  // [23]
    8'd41,  // [24]
    8'd42,  // [25]
    8'd43,  // [26]
    8'd0,   // [27]
    8'd0,   // [28]
    8'd0,   // [29]
    8'd0,   // [30]
    8'd0,   // [31]
    8'd0,   // [32]
    8'd8,   // [33]
    8'd16,  // [34]
    8'd24,  // [35]
    8'd32,  // [36]
    8'd44,  // [37]
    8'd45,  // [38]
    8'd46,  // [39]
    8'd47,  // [40]
    8'd48,  // [41]
    8'd49,  // [42]
    8'd0,   // [43]
    8'd0,   // [44]
    8'd0,   // [45]
    8'd0,   // [46]
    8'd0,   // [47]
    8'd0,   // [48]
    8'd9,   // [49]
    8'd19,  // [50]
    8'd33,  // [51]
    8'd50,  // [52]
    8'd51,  // [53]
    8'd52,  // [54]
    8'd53,  // [55]
    8'd54,  // [56]
    8'd55,  // [57]
    8'd56,  // [58]
    8'd0,   // [59]
    8'd0,   // [60]
    8'd0,   // [61]
    8'd0,   // [62]
    8'd0,   // [63]
    8'd0,   // [64]
    8'd10,  // [65]
    8'd25,  // [66]
    8'd57,  // [67]
    8'd58,  // [68]
    8'd59,  // [69]
    8'd60,  // [70]
    8'd61,  // [71]
    8'd62,  // [72]
    8'd63,  // [73]
    8'd64,  // [74]
    8'd0,   // [75]
    8'd0,   // [76]
    8'd0,   // [77]
    8'd0,   // [78]
    8'd0,   // [79]
    8'd0,   // [80]
    8'd13,  // [81]
    8'd29,  // [82]
    8'd65,  // [83]
    8'd66,  // [84]
    8'd67,  // [85]
    8'd68,  // [86]
    8'd69,  // [87]
    8'd70,  // [88]
    8'd71,  // [89]
    8'd72,  // [90]
    8'd0,   // [91]
    8'd0,   // [92]
    8'd0,   // [93]
    8'd0,   // [94]
    8'd0,   // [95]
    8'd0,   // [96]
    8'd14,  // [97]
    8'd34,  // [98]
    8'd73,  // [99]
    8'd74,  // [100]
    8'd75,  // [101]
    8'd76,  // [102]
    8'd77,  // [103]
    8'd78,  // [104]
    8'd79,  // [105]
    8'd80,  // [106]
    8'd0,   // [107]
    8'd0,   // [108]
    8'd0,   // [109]
    8'd0,   // [110]
    8'd0,   // [111]
    8'd0,   // [112]
    8'd17,  // [113]
    8'd35,  // [114]
    8'd81,  // [115]
    8'd82,  // [116]
    8'd83,  // [117]
    8'd84,  // [118]
    8'd85,  // [119]
    8'd86,  // [120]
    8'd87,  // [121]
    8'd88,  // [122]
    8'd0,   // [123]
    8'd0,   // [124]
    8'd0,   // [125]
    8'd0,   // [126]
    8'd0,   // [127]
    8'd0,   // [128]
    8'd20,  // [129]
    8'd36,  // [130]
    8'd89,  // [131]
    8'd90,  // [132]
    8'd91,  // [133]
    8'd92,  // [134]
    8'd93,  // [135]
    8'd94,  // [136]
    8'd95,  // [137]
    8'd96,  // [138]
    8'd0,   // [139]
    8'd0,   // [140]
    8'd0,   // [141]
    8'd0,   // [142]
    8'd0,   // [143]
    8'd0,   // [144]
    8'd21,  // [145]
    8'd97,  // [146]
    8'd98,  // [147]
    8'd99,  // [148]
    8'd100, // [149]
    8'd101, // [150]
    8'd102, // [151]
    8'd103, // [152]
    8'd104, // [153]
    8'd105, // [154]
    8'd0,   // [155]
    8'd0,   // [156]
    8'd0,   // [157]
    8'd0,   // [158]
    8'd0,   // [159]
    8'd0,   // [160]
    8'd22,  // [161]
    8'd106, // [162]
    8'd107, // [163]
    8'd108, // [164]
    8'd109, // [165]
    8'd110, // [166]
    8'd111, // [167]
    8'd112, // [168]
    8'd113, // [169]
    8'd114, // [170]
    8'd0,   // [171]
    8'd0,   // [172]
    8'd0,   // [173]
    8'd0,   // [174]
    8'd0,   // [175]
    8'd0,   // [176]
    8'd26,  // [177]
    8'd115, // [178]
    8'd116, // [179]
    8'd117, // [180]
    8'd118, // [181]
    8'd119, // [182]
    8'd120, // [183]
    8'd121, // [184]
    8'd122, // [185]
    8'd123, // [186]
    8'd0,   // [187]
    8'd0,   // [188]
    8'd0,   // [189]
    8'd0,   // [190]
    8'd0,   // [191]
    8'd0,   // [192]
    8'd27,  // [193]
    8'd124, // [194]
    8'd125, // [195]
    8'd126, // [196]
    8'd127, // [197]
    8'd128, // [198]
    8'd129, // [199]
    8'd130, // [200]
    8'd131, // [201]
    8'd132, // [202]
    8'd0,   // [203]
    8'd0,   // [204]
    8'd0,   // [205]
    8'd0,   // [206]
    8'd0,   // [207]
    8'd0,   // [208]
    8'd30,  // [209]
    8'd133, // [210]
    8'd134, // [211]
    8'd135, // [212]
    8'd136, // [213]
    8'd137, // [214]
    8'd138, // [215]
    8'd139, // [216]
    8'd140, // [217]
    8'd141, // [218]
    8'd0,   // [219]
    8'd0,   // [220]
    8'd0,   // [221]
    8'd0,   // [222]
    8'd0,   // [223]
    8'd0,   // [224]
    8'd142, // [225]
    8'd143, // [226]
    8'd144, // [227]
    8'd145, // [228]
    8'd146, // [229]
    8'd147, // [230]
    8'd148, // [231]
    8'd149, // [232]
    8'd150, // [233]
    8'd151, // [234]
    8'd0,   // [235]
    8'd0,   // [236]
    8'd0,   // [237]
    8'd0,   // [238]
    8'd0,   // [239]
    8'd31,  // [240]
    8'd152, // [241]
    8'd153, // [242]
    8'd154, // [243]
    8'd155, // [244]
    8'd156, // [245]
    8'd157, // [246]
    8'd158, // [247]
    8'd159, // [248]
    8'd160, // [249]
    8'd161  // [250]
};

`endif //Cb_ HUFF_CONSTANTS_SVH
