`timescale 1ps/1ps

module jpeg_top_TB;

    // ----------------------
    // Declarations
    // ----------------------
    logic end_of_file_signal;
    logic [23:0] data_in;
    logic clk;
    logic rst;
    logic enable;
  logic bitstream_completed;
    wire [31:0] JPEG_bitstream;
    wire data_ready;
    wire [4:0] end_of_file_bitstream_count;
    wire eof_data_partial_ready;

    integer outfile;

    // ----------------------
    // Unit Under Test
    // ----------------------
    jpeg_top UUT (
        .end_of_file_signal(end_of_file_signal),
        .data_in(data_in),
        .clk(clk),
        .rst(rst),
        .enable(enable),
        .JPEG_bitstream(JPEG_bitstream),
        .data_ready(data_ready),
        .end_of_file_bitstream_count(end_of_file_bitstream_count),
        .eof_data_partial_ready(eof_data_partial_ready)
    );

    // ----------------------
    // Stimulus process
    // ----------------------
    initial begin : STIMUL
        rst = 1'b1;
        enable = 1'b0;
        end_of_file_signal = 1'b0;
        data_in = '0;
   bitstream_completed = 1'b0;
        #10000;
        rst = 1'b0;
        enable = 1'b1;

 // Insert pixel data generated by Python

     `include "pixel_data.txt"



        #130000;
        enable = 1'b0;
        #2000000;
	     bitstream_completed = 1'b1;
    end

    // ----------------------
    // Open output file once
    // ----------------------
    initial begin

       outfile = $fopen("raw_jpeg_bitstream_to_image/bitstream_output.txt", "w");
        if (outfile == 0) begin
            $display("ERROR: Could not open bitstream_output.txt");
            $finish;
        end
    end

    // ----------------------
    // End simulation when JPEG bitstream = 0
    // ----------------------
    always_ff @(posedge clk) begin
        if (data_ready) begin
            if (   bitstream_completed == 1'b1) begin
                $display("INFO: End of JPEG stream detected. Closing file and stopping.");
                $fclose(outfile);
                $finish;
            end
        end
    end

    // ----------------------
    // Clock generator
    // ----------------------
    always begin : CLOCK_clk
        clk = 1'b0;
        #5000;
        clk = 1'b1;
        #5000;
    end

    // ----------------------
    // Write JPEG bitstream whenever ready
    // ----------------------
    always_ff @(posedge clk) begin : JPEG
        if (data_ready) begin
            $fwrite(outfile, "%h\n", JPEG_bitstream);   // write in hex
        end
    end

endmodule
