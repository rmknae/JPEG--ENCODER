// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
//    Header file defining localparams for JPEG Huffman encoding.
//    - DC Huffman code lengths and codes (Luma & Chroma)
//    - AC Huffman code lengths and codes (Luma & Chroma)
//    - Run-length/size to Huffman index mapping
//
// Author: Rameen
// Date  : 23rd July 2025

`ifndef HUFF_CONSTANTS_SVH
`define HUFF_CONSTANTS_SVH


`endif // HUFF_CONSTANTS_SVH
