// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
//    Header file defining localparams for JPEG Huffman encoding.
//    - DC Huffman code lengths and codes (Luma & Chroma)
//    - AC Huffman code lengths and codes (Luma & Chroma)
//    - Run-length/size to Huffman index mapping
//
// Author: Rameen
// Date  : 23rd July 2025

`ifndef Y_HUFF_CONSTANTS_SVH
`define Y_HUFF_CONSTANTS_SVH
// ====================================================================
// Y Component Huffman Table Constants
// Automatically generated from JPEG Huffman tables
// Include this file in your module with: `include "y_huffman_constants.svh`
// ====================================================================

// -------------------- DC Code Lengths --------------------
parameter int Y_DC_code_length[0:11] = '{2,2,2,3,4,5,6,7,8,9,10,11};

// -------------------- DC Codes --------------------
parameter logic [10:0] Y_DC[0:11] = '{
    11'b00000000000, 11'b01000000000, 11'b10000000000, 11'b11000000000,
    11'b11100000000, 11'b11110000000, 11'b11111000000, 11'b11111100000,
    11'b11111110000, 11'b11111111000, 11'b11111111100, 11'b11111111110
};

// -------------------- AC Code Lengths --------------------
parameter int Y_AC_code_length[0:161] = '{
    2,2,3,4,4,4,5,5,5,6,6,7,7,7,7,8,
    8,8,9,9,9,9,9,10,10,10,10,10,11,11,11,11,
    12,12,12,12,15,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,
    16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16
};

// -------------------- AC Codes --------------------
parameter logic [15:0] Y_AC[0:161] = '{
    16'b0000000000000000, 16'b0100000000000000, 16'b1000000000000000, 16'b1010000000000000,
    16'b1011000000000000, 16'b1100000000000000, 16'b1101000000000000, 16'b1101100000000000,
    16'b1110000000000000, 16'b1110100000000000, 16'b1110110000000000, 16'b1111000000000000,
    16'b1111001000000000, 16'b1111010000000000, 16'b1111011000000000, 16'b1111100000000000,
    16'b1111100100000000, 16'b1111101000000000, 16'b1111101100000000, 16'b1111101110000000,
    16'b1111110000000000, 16'b1111110010000000, 16'b1111110100000000, 16'b1111110110000000,
    16'b1111110111000000, 16'b1111111000000000, 16'b1111111001000000, 16'b1111111010000000,
    16'b1111111011000000, 16'b1111111011100000, 16'b1111111100000000, 16'b1111111100100000,
    16'b1111111101000000, 16'b1111111101010000, 16'b1111111101100000, 16'b1111111101110000,
    16'b1111111110000000, 16'b1111111110000010, 16'b1111111110000011, 16'b1111111110000100,
    16'b1111111110000101, 16'b1111111110000110, 16'b1111111110000111, 16'b1111111110001000,
    16'b1111111110001001, 16'b1111111110001010, 16'b1111111110001011, 16'b1111111110001100,
    16'b1111111110001101, 16'b1111111110001110, 16'b1111111110001111, 16'b1111111110010000,
    16'b1111111110010001, 16'b1111111110010010, 16'b1111111110010011, 16'b1111111110010100,
    16'b1111111110010101, 16'b1111111110010110, 16'b1111111110010111, 16'b1111111110011000,
    16'b1111111110011001, 16'b1111111110011010, 16'b1111111110011011, 16'b1111111110011100,
    16'b1111111110011101, 16'b1111111110011110, 16'b1111111110011111, 16'b1111111110100000,
    16'b1111111110100001, 16'b1111111110100010, 16'b1111111110100011, 16'b1111111110100100,
    16'b1111111110100101, 16'b1111111110100110, 16'b1111111110100111, 16'b1111111110101000,
    16'b1111111110101001, 16'b1111111110101010, 16'b1111111110101011, 16'b1111111110101100,
    16'b1111111110101101, 16'b1111111110101110, 16'b1111111110101111, 16'b1111111110110000,
    16'b1111111110110001, 16'b1111111110110010, 16'b1111111110110011, 16'b1111111110110100,
    16'b1111111110110101, 16'b1111111110110110, 16'b1111111110110111, 16'b1111111110111000,
    16'b1111111110111001, 16'b1111111110111010, 16'b1111111110111011, 16'b1111111110111100,
    16'b1111111110111101, 16'b1111111110111110, 16'b1111111110111111, 16'b1111111111000000,
    16'b1111111111000001, 16'b1111111111000010, 16'b1111111111000011, 16'b1111111111000100,
    16'b1111111111000101, 16'b1111111111000110, 16'b1111111111000111, 16'b1111111111001000,
    16'b1111111111001001, 16'b1111111111001010, 16'b1111111111001011, 16'b1111111111001100,
    16'b1111111111001101, 16'b1111111111001110, 16'b1111111111001111, 16'b1111111111010000,
    16'b1111111111010001, 16'b1111111111010010, 16'b1111111111010011, 16'b1111111111010100,
    16'b1111111111010101, 16'b1111111111010110, 16'b1111111111010111, 16'b1111111111011000,
    16'b1111111111011001, 16'b1111111111011010, 16'b1111111111011011, 16'b1111111111011100,
    16'b1111111111011101, 16'b1111111111011110, 16'b1111111111011111, 16'b1111111111100000,
    16'b1111111111100001, 16'b1111111111100010, 16'b1111111111100011, 16'b1111111111100100,
    16'b1111111111100101, 16'b1111111111100110, 16'b1111111111100111, 16'b1111111111101000,
    16'b1111111111101001, 16'b1111111111101010, 16'b1111111111101011, 16'b1111111111101100,
    16'b1111111111101101, 16'b1111111111101110, 16'b1111111111101111, 16'b1111111111110000,
    16'b1111111111110001, 16'b1111111111110010, 16'b1111111111110011, 16'b1111111111110100,
    16'b1111111111110101, 16'b1111111111110110, 16'b1111111111110111, 16'b1111111111111000,
    16'b1111111111111001, 16'b1111111111111010, 16'b1111111111111011, 16'b1111111111111100,
    16'b1111111111111101, 16'b1111111111111110
};



`endif //y_ HUFF_CONSTANTS_SVH
