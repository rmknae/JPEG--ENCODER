// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file // for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
//   Defines the standard JPEG luminance quantization matrix (8x8)  //  used for testing quantizer modules.
//
// Author : Navaal Noshi
// Date   : 29th July 2025
//

`ifndef QUANTIZER_CONSTANTS_SVH
`define QUANTIZER_CONSTANTS_SVH



`endif // QUANTIZER_CONSTANTS_SVH
